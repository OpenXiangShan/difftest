module AXI4FakeDMA(
  input          clock,
  input          reset,
  input          auto_dma_out_awready,
  output         auto_dma_out_awvalid,
  output [7:0]   auto_dma_out_awid,
  output [37:0]  auto_dma_out_awaddr,
  input          auto_dma_out_wready,
  output         auto_dma_out_wvalid,
  output [255:0] auto_dma_out_wdata,
  output [31:0]  auto_dma_out_wstrb,
  output         auto_dma_out_wlast,
  input          auto_dma_out_bvalid,
  input  [7:0]   auto_dma_out_bid,
  input          auto_dma_out_arready,
  output         auto_dma_out_arvalid,
  output [7:0]   auto_dma_out_arid,
  output [37:0]  auto_dma_out_araddr,
  input          auto_dma_out_rvalid,
  input  [7:0]   auto_dma_out_rid,
  input  [255:0] auto_dma_out_rdata,
  output         auto_in_awready,
  input          auto_in_awvalid,
  input          auto_in_awid,
  input  [36:0]  auto_in_awaddr,
  input  [7:0]   auto_in_awlen,
  input  [2:0]   auto_in_awsize,
  input  [1:0]   auto_in_awburst,
  input          auto_in_awlock,
  input  [3:0]   auto_in_awcache,
  input  [2:0]   auto_in_awprot,
  input  [3:0]   auto_in_awqos,
  output         auto_in_wready,
  input          auto_in_wvalid,
  input  [63:0]  auto_in_wdata,
  input  [7:0]   auto_in_wstrb,
  input          auto_in_wlast,
  input          auto_in_bready,
  output         auto_in_bvalid,
  output         auto_in_bid,
  output [1:0]   auto_in_bresp,
  output         auto_in_arready,
  input          auto_in_arvalid,
  input          auto_in_arid,
  input  [36:0]  auto_in_araddr,
  input  [7:0]   auto_in_arlen,
  input  [2:0]   auto_in_arsize,
  input  [1:0]   auto_in_arburst,
  input          auto_in_arlock,
  input  [3:0]   auto_in_arcache,
  input  [2:0]   auto_in_arprot,
  input  [3:0]   auto_in_arqos,
  input          auto_in_rready,
  output         auto_in_rvalid,
  output         auto_in_rid,
  output [63:0]  auto_in_rdata,
  output [1:0]   auto_in_rresp,
  output         auto_in_rlast
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [511:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  wire  mshr_0_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_0_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_0_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_0_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_0_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_0_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_0_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_0_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_0_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_0_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_0_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_0_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_0_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_0_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_0_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_1_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_1_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_1_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_1_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_1_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_1_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_1_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_1_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_1_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_1_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_1_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_1_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_1_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_1_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_1_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_2_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_2_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_2_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_2_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_2_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_2_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_2_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_2_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_2_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_2_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_2_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_2_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_2_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_2_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_2_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_3_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_3_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_3_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_3_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_3_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_3_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_3_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_3_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_3_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_3_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_3_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_3_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_3_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_3_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_3_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_4_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_4_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_4_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_4_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_4_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_4_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_4_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_4_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_4_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_4_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_4_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_4_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_4_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_4_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_4_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_5_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_5_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_5_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_5_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_5_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_5_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_5_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_5_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_5_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_5_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_5_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_5_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_5_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_5_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_5_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_6_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_6_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_6_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_6_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_6_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_6_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_6_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_6_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_6_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_6_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_6_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_6_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_6_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_6_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_6_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_7_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_7_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_7_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_7_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_7_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_7_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_7_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_7_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_7_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_7_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_7_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_7_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_7_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_7_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_7_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_8_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_8_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_8_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_8_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_8_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_8_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_8_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_8_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_8_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_8_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_8_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_8_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_8_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_8_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_8_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_9_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_9_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_9_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_9_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_9_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_9_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_9_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_9_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_9_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_9_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_9_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_9_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_9_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_9_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_9_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_10_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_10_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_10_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_10_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_10_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_10_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_10_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_10_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_10_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_10_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_10_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_10_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_10_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_10_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_10_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_11_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_11_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_11_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_11_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_11_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_11_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_11_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_11_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_11_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_11_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_11_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_11_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_11_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_11_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_11_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_12_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_12_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_12_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_12_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_12_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_12_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_12_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_12_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_12_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_12_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_12_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_12_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_12_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_12_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_12_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_13_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_13_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_13_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_13_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_13_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_13_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_13_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_13_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_13_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_13_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_13_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_13_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_13_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_13_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_13_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_14_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_14_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_14_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_14_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_14_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_14_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_14_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_14_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_14_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_14_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_14_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_14_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_14_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_14_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_14_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_15_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_15_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_15_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_15_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_15_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_15_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_15_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_15_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_15_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_15_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_15_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_15_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_15_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_15_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_15_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_16_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_16_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_16_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_16_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_16_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_16_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_16_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_16_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_16_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_16_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_16_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_16_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_16_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_16_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_16_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_17_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_17_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_17_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_17_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_17_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_17_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_17_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_17_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_17_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_17_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_17_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_17_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_17_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_17_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_17_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_18_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_18_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_18_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_18_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_18_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_18_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_18_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_18_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_18_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_18_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_18_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_18_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_18_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_18_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_18_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_19_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_19_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_19_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_19_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_19_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_19_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_19_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_19_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_19_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_19_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_19_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_19_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_19_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_19_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_19_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_20_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_20_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_20_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_20_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_20_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_20_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_20_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_20_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_20_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_20_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_20_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_20_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_20_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_20_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_20_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_21_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_21_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_21_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_21_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_21_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_21_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_21_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_21_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_21_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_21_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_21_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_21_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_21_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_21_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_21_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_22_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_22_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_22_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_22_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_22_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_22_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_22_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_22_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_22_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_22_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_22_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_22_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_22_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_22_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_22_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_23_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_23_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_23_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_23_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_23_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_23_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_23_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_23_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_23_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_23_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_23_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_23_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_23_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_23_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_23_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_24_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_24_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_24_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_24_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_24_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_24_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_24_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_24_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_24_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_24_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_24_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_24_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_24_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_24_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_24_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_25_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_25_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_25_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_25_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_25_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_25_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_25_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_25_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_25_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_25_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_25_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_25_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_25_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_25_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_25_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_26_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_26_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_26_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_26_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_26_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_26_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_26_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_26_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_26_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_26_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_26_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_26_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_26_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_26_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_26_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_27_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_27_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_27_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_27_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_27_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_27_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_27_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_27_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_27_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_27_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_27_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_27_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_27_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_27_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_27_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_28_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_28_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_28_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_28_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_28_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_28_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_28_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_28_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_28_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_28_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_28_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_28_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_28_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_28_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_28_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_29_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_29_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_29_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_29_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_29_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_29_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_29_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_29_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_29_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_29_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_29_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_29_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_29_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_29_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_29_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_30_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_30_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_30_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_30_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_30_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_30_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_30_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_30_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_30_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_30_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_30_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_30_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_30_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_30_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_30_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_31_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_31_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_31_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_31_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_31_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_31_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_31_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_31_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_31_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_31_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_31_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_31_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_31_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_31_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_31_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_32_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_32_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_32_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_32_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_32_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_32_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_32_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_32_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_32_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_32_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_32_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_32_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_32_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_32_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_32_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_33_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_33_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_33_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_33_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_33_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_33_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_33_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_33_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_33_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_33_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_33_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_33_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_33_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_33_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_33_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_34_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_34_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_34_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_34_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_34_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_34_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_34_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_34_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_34_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_34_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_34_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_34_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_34_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_34_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_34_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_35_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_35_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_35_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_35_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_35_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_35_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_35_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_35_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_35_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_35_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_35_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_35_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_35_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_35_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_35_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_36_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_36_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_36_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_36_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_36_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_36_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_36_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_36_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_36_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_36_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_36_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_36_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_36_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_36_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_36_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_37_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_37_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_37_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_37_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_37_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_37_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_37_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_37_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_37_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_37_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_37_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_37_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_37_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_37_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_37_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_38_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_38_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_38_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_38_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_38_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_38_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_38_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_38_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_38_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_38_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_38_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_38_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_38_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_38_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_38_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_39_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_39_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_39_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_39_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_39_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_39_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_39_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_39_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_39_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_39_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_39_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_39_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_39_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_39_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_39_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_40_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_40_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_40_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_40_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_40_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_40_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_40_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_40_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_40_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_40_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_40_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_40_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_40_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_40_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_40_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_41_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_41_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_41_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_41_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_41_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_41_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_41_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_41_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_41_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_41_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_41_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_41_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_41_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_41_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_41_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_42_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_42_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_42_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_42_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_42_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_42_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_42_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_42_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_42_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_42_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_42_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_42_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_42_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_42_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_42_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_43_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_43_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_43_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_43_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_43_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_43_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_43_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_43_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_43_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_43_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_43_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_43_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_43_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_43_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_43_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_44_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_44_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_44_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_44_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_44_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_44_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_44_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_44_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_44_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_44_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_44_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_44_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_44_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_44_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_44_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_45_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_45_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_45_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_45_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_45_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_45_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_45_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_45_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_45_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_45_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_45_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_45_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_45_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_45_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_45_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_46_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_46_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_46_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_46_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_46_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_46_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_46_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_46_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_46_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_46_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_46_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_46_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_46_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_46_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_46_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_47_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_47_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_47_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_47_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_47_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_47_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_47_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_47_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_47_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_47_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_47_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_47_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_47_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_47_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_47_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_48_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_48_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_48_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_48_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_48_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_48_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_48_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_48_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_48_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_48_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_48_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_48_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_48_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_48_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_48_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_49_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_49_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_49_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_49_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_49_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_49_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_49_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_49_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_49_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_49_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_49_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_49_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_49_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_49_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_49_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_50_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_50_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_50_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_50_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_50_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_50_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_50_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_50_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_50_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_50_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_50_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_50_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_50_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_50_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_50_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_51_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_51_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_51_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_51_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_51_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_51_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_51_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_51_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_51_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_51_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_51_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_51_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_51_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_51_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_51_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_52_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_52_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_52_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_52_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_52_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_52_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_52_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_52_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_52_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_52_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_52_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_52_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_52_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_52_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_52_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_53_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_53_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_53_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_53_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_53_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_53_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_53_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_53_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_53_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_53_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_53_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_53_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_53_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_53_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_53_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_54_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_54_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_54_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_54_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_54_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_54_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_54_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_54_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_54_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_54_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_54_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_54_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_54_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_54_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_54_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_55_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_55_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_55_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_55_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_55_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_55_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_55_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_55_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_55_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_55_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_55_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_55_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_55_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_55_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_55_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_56_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_56_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_56_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_56_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_56_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_56_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_56_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_56_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_56_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_56_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_56_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_56_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_56_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_56_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_56_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_57_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_57_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_57_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_57_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_57_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_57_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_57_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_57_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_57_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_57_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_57_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_57_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_57_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_57_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_57_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_58_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_58_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_58_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_58_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_58_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_58_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_58_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_58_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_58_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_58_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_58_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_58_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_58_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_58_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_58_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_59_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_59_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_59_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_59_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_59_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_59_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_59_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_59_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_59_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_59_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_59_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_59_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_59_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_59_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_59_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_60_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_60_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_60_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_60_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_60_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_60_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_60_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_60_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_60_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_60_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_60_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_60_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_60_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_60_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_60_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_61_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_61_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_61_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_61_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_61_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_61_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_61_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_61_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_61_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_61_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_61_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_61_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_61_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_61_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_61_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_62_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_62_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_62_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_62_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_62_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_62_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_62_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_62_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_62_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_62_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_62_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_62_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_62_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_62_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_62_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_63_clock; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_63_reset; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_63_io_enable; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_63_io_slave_wen; // @[AXI4FakeDMA.scala 149:44]
  wire [3:0] mshr_63_io_slave_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_63_io_slave_rdata; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_63_io_slave_wdata; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_63_io_master_req_valid; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_63_io_master_req_ready; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_63_io_master_req_is_write; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_63_io_master_req_addr; // @[AXI4FakeDMA.scala 149:44]
  wire [63:0] mshr_63_io_master_req_mask; // @[AXI4FakeDMA.scala 149:44]
  wire [511:0] mshr_63_io_master_req_data; // @[AXI4FakeDMA.scala 149:44]
  wire  mshr_63_io_master_resp_valid; // @[AXI4FakeDMA.scala 149:44]
  wire [255:0] mshr_63_io_master_resp_bits; // @[AXI4FakeDMA.scala 149:44]
  reg [1:0] state; // @[AXI4SlaveModule.scala 95:22]
  wire  _bundleIn_0_arready_T = state == 2'h0; // @[AXI4SlaveModule.scala 153:24]
  wire  in_arready = state == 2'h0; // @[AXI4SlaveModule.scala 153:24]
  wire  in_arvalid = auto_in_arvalid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  wire  _T = in_arready & in_arvalid; // @[Decoupled.scala 50:35]
  wire  in_awready = _bundleIn_0_arready_T & ~in_arvalid; // @[AXI4SlaveModule.scala 171:35]
  wire  in_awvalid = auto_in_awvalid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  wire  _T_1 = in_awready & in_awvalid; // @[Decoupled.scala 50:35]
  wire  in_wready = state == 2'h2; // @[AXI4SlaveModule.scala 172:23]
  wire  in_wvalid = auto_in_wvalid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  wire  _T_2 = in_wready & in_wvalid; // @[Decoupled.scala 50:35]
  wire  in_bready = auto_in_bready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  wire  in_bvalid = state == 2'h3; // @[AXI4SlaveModule.scala 175:22]
  wire  _T_3 = in_bready & in_bvalid; // @[Decoupled.scala 50:35]
  wire  in_rready = auto_in_rready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  wire  in_rvalid = state == 2'h1; // @[AXI4SlaveModule.scala 155:23]
  wire  _T_4 = in_rready & in_rvalid; // @[Decoupled.scala 50:35]
  wire [1:0] in_awburst = auto_in_awburst; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  wire [1:0] in_arburst = auto_in_arburst; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  reg [7:0] value; // @[Counter.scala 62:40]
  wire [7:0] in_arlen = auto_in_arlen; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  reg [7:0] hold_data; // @[Reg.scala 16:16]
  wire [7:0] _T_27 = _T ? in_arlen : hold_data; // @[Hold.scala 25:8]
  wire  in_rlast = value == _T_27; // @[AXI4SlaveModule.scala 133:32]
  wire  in_wlast = auto_in_wlast; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  wire [1:0] _GEN_3 = _T_2 & in_wlast ? 2'h3 : state; // @[AXI4SlaveModule.scala 112:42 113:15 95:22]
  wire [1:0] _GEN_4 = _T_3 ? 2'h0 : state; // @[AXI4SlaveModule.scala 117:24 118:15 95:22]
  wire [1:0] _GEN_5 = 2'h3 == state ? _GEN_4 : state; // @[AXI4SlaveModule.scala 97:16 95:22]
  wire [7:0] in_wstrb = auto_in_wstrb; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  reg [36:0] raddr_hold_data; // @[Reg.scala 16:16]
  wire [36:0] in_araddr = auto_in_araddr; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  wire [36:0] _GEN_10 = _T ? in_araddr : raddr_hold_data; // @[Reg.scala 16:16 17:{18,22}]
  wire [7:0] _value_T_1 = value + 8'h1; // @[Counter.scala 78:24]
  reg [36:0] waddr_hold_data; // @[Reg.scala 16:16]
  wire [36:0] in_awaddr = auto_in_awaddr; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  wire [36:0] _GEN_13 = _T_1 ? in_awaddr : waddr_hold_data; // @[Reg.scala 16:16 17:{18,22}]
  reg  bundleIn_0_bid_r; // @[Reg.scala 16:16]
  wire  in_awid = auto_in_awid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  reg  bundleIn_0_rid_r; // @[Reg.scala 16:16]
  wire  in_arid = auto_in_arid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  reg [63:0] enable; // @[AXI4FakeDMA.scala 151:25]
  wire [3:0] reqReadOffset = _GEN_10[6:3]; // @[AXI4FakeDMA.scala 155:30]
  wire [6:0] reqReadIdx = _GEN_10[13:7]; // @[AXI4FakeDMA.scala 156:27]
  wire [63:0] req_r0 = mshr_0_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] req_r1 = mshr_1_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_19 = 6'h1 == reqReadIdx[5:0] ? req_r1 : req_r0; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r2 = mshr_2_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_20 = 6'h2 == reqReadIdx[5:0] ? req_r2 : _GEN_19; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r3 = mshr_3_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_21 = 6'h3 == reqReadIdx[5:0] ? req_r3 : _GEN_20; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r4 = mshr_4_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_22 = 6'h4 == reqReadIdx[5:0] ? req_r4 : _GEN_21; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r5 = mshr_5_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_23 = 6'h5 == reqReadIdx[5:0] ? req_r5 : _GEN_22; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r6 = mshr_6_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_24 = 6'h6 == reqReadIdx[5:0] ? req_r6 : _GEN_23; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r7 = mshr_7_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_25 = 6'h7 == reqReadIdx[5:0] ? req_r7 : _GEN_24; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r8 = mshr_8_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_26 = 6'h8 == reqReadIdx[5:0] ? req_r8 : _GEN_25; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r9 = mshr_9_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_27 = 6'h9 == reqReadIdx[5:0] ? req_r9 : _GEN_26; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r10 = mshr_10_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_28 = 6'ha == reqReadIdx[5:0] ? req_r10 : _GEN_27; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r11 = mshr_11_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_29 = 6'hb == reqReadIdx[5:0] ? req_r11 : _GEN_28; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r12 = mshr_12_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_30 = 6'hc == reqReadIdx[5:0] ? req_r12 : _GEN_29; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r13 = mshr_13_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_31 = 6'hd == reqReadIdx[5:0] ? req_r13 : _GEN_30; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r14 = mshr_14_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_32 = 6'he == reqReadIdx[5:0] ? req_r14 : _GEN_31; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r15 = mshr_15_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_33 = 6'hf == reqReadIdx[5:0] ? req_r15 : _GEN_32; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r16 = mshr_16_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_34 = 6'h10 == reqReadIdx[5:0] ? req_r16 : _GEN_33; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r17 = mshr_17_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_35 = 6'h11 == reqReadIdx[5:0] ? req_r17 : _GEN_34; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r18 = mshr_18_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_36 = 6'h12 == reqReadIdx[5:0] ? req_r18 : _GEN_35; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r19 = mshr_19_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_37 = 6'h13 == reqReadIdx[5:0] ? req_r19 : _GEN_36; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r20 = mshr_20_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_38 = 6'h14 == reqReadIdx[5:0] ? req_r20 : _GEN_37; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r21 = mshr_21_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_39 = 6'h15 == reqReadIdx[5:0] ? req_r21 : _GEN_38; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r22 = mshr_22_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_40 = 6'h16 == reqReadIdx[5:0] ? req_r22 : _GEN_39; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r23 = mshr_23_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_41 = 6'h17 == reqReadIdx[5:0] ? req_r23 : _GEN_40; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r24 = mshr_24_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_42 = 6'h18 == reqReadIdx[5:0] ? req_r24 : _GEN_41; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r25 = mshr_25_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_43 = 6'h19 == reqReadIdx[5:0] ? req_r25 : _GEN_42; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r26 = mshr_26_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_44 = 6'h1a == reqReadIdx[5:0] ? req_r26 : _GEN_43; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r27 = mshr_27_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_45 = 6'h1b == reqReadIdx[5:0] ? req_r27 : _GEN_44; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r28 = mshr_28_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_46 = 6'h1c == reqReadIdx[5:0] ? req_r28 : _GEN_45; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r29 = mshr_29_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_47 = 6'h1d == reqReadIdx[5:0] ? req_r29 : _GEN_46; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r30 = mshr_30_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_48 = 6'h1e == reqReadIdx[5:0] ? req_r30 : _GEN_47; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r31 = mshr_31_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_49 = 6'h1f == reqReadIdx[5:0] ? req_r31 : _GEN_48; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r32 = mshr_32_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_50 = 6'h20 == reqReadIdx[5:0] ? req_r32 : _GEN_49; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r33 = mshr_33_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_51 = 6'h21 == reqReadIdx[5:0] ? req_r33 : _GEN_50; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r34 = mshr_34_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_52 = 6'h22 == reqReadIdx[5:0] ? req_r34 : _GEN_51; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r35 = mshr_35_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_53 = 6'h23 == reqReadIdx[5:0] ? req_r35 : _GEN_52; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r36 = mshr_36_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_54 = 6'h24 == reqReadIdx[5:0] ? req_r36 : _GEN_53; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r37 = mshr_37_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_55 = 6'h25 == reqReadIdx[5:0] ? req_r37 : _GEN_54; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r38 = mshr_38_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_56 = 6'h26 == reqReadIdx[5:0] ? req_r38 : _GEN_55; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r39 = mshr_39_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_57 = 6'h27 == reqReadIdx[5:0] ? req_r39 : _GEN_56; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r40 = mshr_40_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_58 = 6'h28 == reqReadIdx[5:0] ? req_r40 : _GEN_57; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r41 = mshr_41_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_59 = 6'h29 == reqReadIdx[5:0] ? req_r41 : _GEN_58; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r42 = mshr_42_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_60 = 6'h2a == reqReadIdx[5:0] ? req_r42 : _GEN_59; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r43 = mshr_43_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_61 = 6'h2b == reqReadIdx[5:0] ? req_r43 : _GEN_60; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r44 = mshr_44_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_62 = 6'h2c == reqReadIdx[5:0] ? req_r44 : _GEN_61; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r45 = mshr_45_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_63 = 6'h2d == reqReadIdx[5:0] ? req_r45 : _GEN_62; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r46 = mshr_46_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_64 = 6'h2e == reqReadIdx[5:0] ? req_r46 : _GEN_63; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r47 = mshr_47_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_65 = 6'h2f == reqReadIdx[5:0] ? req_r47 : _GEN_64; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r48 = mshr_48_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_66 = 6'h30 == reqReadIdx[5:0] ? req_r48 : _GEN_65; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r49 = mshr_49_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_67 = 6'h31 == reqReadIdx[5:0] ? req_r49 : _GEN_66; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r50 = mshr_50_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_68 = 6'h32 == reqReadIdx[5:0] ? req_r50 : _GEN_67; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r51 = mshr_51_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_69 = 6'h33 == reqReadIdx[5:0] ? req_r51 : _GEN_68; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r52 = mshr_52_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_70 = 6'h34 == reqReadIdx[5:0] ? req_r52 : _GEN_69; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r53 = mshr_53_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_71 = 6'h35 == reqReadIdx[5:0] ? req_r53 : _GEN_70; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r54 = mshr_54_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_72 = 6'h36 == reqReadIdx[5:0] ? req_r54 : _GEN_71; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r55 = mshr_55_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_73 = 6'h37 == reqReadIdx[5:0] ? req_r55 : _GEN_72; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r56 = mshr_56_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_74 = 6'h38 == reqReadIdx[5:0] ? req_r56 : _GEN_73; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r57 = mshr_57_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_75 = 6'h39 == reqReadIdx[5:0] ? req_r57 : _GEN_74; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r58 = mshr_58_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_76 = 6'h3a == reqReadIdx[5:0] ? req_r58 : _GEN_75; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r59 = mshr_59_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_77 = 6'h3b == reqReadIdx[5:0] ? req_r59 : _GEN_76; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r60 = mshr_60_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_78 = 6'h3c == reqReadIdx[5:0] ? req_r60 : _GEN_77; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r61 = mshr_61_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_79 = 6'h3d == reqReadIdx[5:0] ? req_r61 : _GEN_78; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r62 = mshr_62_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_80 = 6'h3e == reqReadIdx[5:0] ? req_r62 : _GEN_79; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [63:0] req_r63 = mshr_63_io_slave_rdata; // @[AXI4FakeDMA.scala 157:{24,24}]
  wire [63:0] _GEN_81 = 6'h3f == reqReadIdx[5:0] ? req_r63 : _GEN_80; // @[AXI4FakeDMA.scala 158:{26,26}]
  wire [3:0] reqWriteOffset = _GEN_13[6:3]; // @[AXI4FakeDMA.scala 161:31]
  wire [6:0] reqWriteIdx = _GEN_13[13:7]; // @[AXI4FakeDMA.scala 162:28]
  wire [63:0] in_wdata = auto_in_wdata; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  wire  has_read_req_0 = mshr_0_io_master_req_valid & ~mshr_0_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_1 = mshr_1_io_master_req_valid & ~mshr_1_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_2 = mshr_2_io_master_req_valid & ~mshr_2_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_3 = mshr_3_io_master_req_valid & ~mshr_3_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_4 = mshr_4_io_master_req_valid & ~mshr_4_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_5 = mshr_5_io_master_req_valid & ~mshr_5_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_6 = mshr_6_io_master_req_valid & ~mshr_6_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_7 = mshr_7_io_master_req_valid & ~mshr_7_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_8 = mshr_8_io_master_req_valid & ~mshr_8_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_9 = mshr_9_io_master_req_valid & ~mshr_9_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_10 = mshr_10_io_master_req_valid & ~mshr_10_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_11 = mshr_11_io_master_req_valid & ~mshr_11_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_12 = mshr_12_io_master_req_valid & ~mshr_12_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_13 = mshr_13_io_master_req_valid & ~mshr_13_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_14 = mshr_14_io_master_req_valid & ~mshr_14_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_15 = mshr_15_io_master_req_valid & ~mshr_15_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_16 = mshr_16_io_master_req_valid & ~mshr_16_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_17 = mshr_17_io_master_req_valid & ~mshr_17_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_18 = mshr_18_io_master_req_valid & ~mshr_18_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_19 = mshr_19_io_master_req_valid & ~mshr_19_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_20 = mshr_20_io_master_req_valid & ~mshr_20_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_21 = mshr_21_io_master_req_valid & ~mshr_21_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_22 = mshr_22_io_master_req_valid & ~mshr_22_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_23 = mshr_23_io_master_req_valid & ~mshr_23_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_24 = mshr_24_io_master_req_valid & ~mshr_24_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_25 = mshr_25_io_master_req_valid & ~mshr_25_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_26 = mshr_26_io_master_req_valid & ~mshr_26_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_27 = mshr_27_io_master_req_valid & ~mshr_27_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_28 = mshr_28_io_master_req_valid & ~mshr_28_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_29 = mshr_29_io_master_req_valid & ~mshr_29_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_30 = mshr_30_io_master_req_valid & ~mshr_30_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_31 = mshr_31_io_master_req_valid & ~mshr_31_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_32 = mshr_32_io_master_req_valid & ~mshr_32_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_33 = mshr_33_io_master_req_valid & ~mshr_33_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_34 = mshr_34_io_master_req_valid & ~mshr_34_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_35 = mshr_35_io_master_req_valid & ~mshr_35_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_36 = mshr_36_io_master_req_valid & ~mshr_36_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_37 = mshr_37_io_master_req_valid & ~mshr_37_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_38 = mshr_38_io_master_req_valid & ~mshr_38_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_39 = mshr_39_io_master_req_valid & ~mshr_39_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_40 = mshr_40_io_master_req_valid & ~mshr_40_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_41 = mshr_41_io_master_req_valid & ~mshr_41_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_42 = mshr_42_io_master_req_valid & ~mshr_42_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_43 = mshr_43_io_master_req_valid & ~mshr_43_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_44 = mshr_44_io_master_req_valid & ~mshr_44_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_45 = mshr_45_io_master_req_valid & ~mshr_45_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_46 = mshr_46_io_master_req_valid & ~mshr_46_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_47 = mshr_47_io_master_req_valid & ~mshr_47_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_48 = mshr_48_io_master_req_valid & ~mshr_48_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_49 = mshr_49_io_master_req_valid & ~mshr_49_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_50 = mshr_50_io_master_req_valid & ~mshr_50_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_51 = mshr_51_io_master_req_valid & ~mshr_51_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_52 = mshr_52_io_master_req_valid & ~mshr_52_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_53 = mshr_53_io_master_req_valid & ~mshr_53_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_54 = mshr_54_io_master_req_valid & ~mshr_54_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_55 = mshr_55_io_master_req_valid & ~mshr_55_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_56 = mshr_56_io_master_req_valid & ~mshr_56_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_57 = mshr_57_io_master_req_valid & ~mshr_57_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_58 = mshr_58_io_master_req_valid & ~mshr_58_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_59 = mshr_59_io_master_req_valid & ~mshr_59_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_60 = mshr_60_io_master_req_valid & ~mshr_60_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_61 = mshr_61_io_master_req_valid & ~mshr_61_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_62 = mshr_62_io_master_req_valid & ~mshr_62_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire  has_read_req_63 = mshr_63_io_master_req_valid & ~mshr_63_io_master_req_is_write; // @[AXI4FakeDMA.scala 131:48]
  wire [63:0] _out_read_index_enc_T = has_read_req_63 ? 64'h8000000000000000 : 64'h0; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_1 = has_read_req_62 ? 64'h4000000000000000 : _out_read_index_enc_T; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_2 = has_read_req_61 ? 64'h2000000000000000 : _out_read_index_enc_T_1; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_3 = has_read_req_60 ? 64'h1000000000000000 : _out_read_index_enc_T_2; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_4 = has_read_req_59 ? 64'h800000000000000 : _out_read_index_enc_T_3; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_5 = has_read_req_58 ? 64'h400000000000000 : _out_read_index_enc_T_4; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_6 = has_read_req_57 ? 64'h200000000000000 : _out_read_index_enc_T_5; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_7 = has_read_req_56 ? 64'h100000000000000 : _out_read_index_enc_T_6; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_8 = has_read_req_55 ? 64'h80000000000000 : _out_read_index_enc_T_7; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_9 = has_read_req_54 ? 64'h40000000000000 : _out_read_index_enc_T_8; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_10 = has_read_req_53 ? 64'h20000000000000 : _out_read_index_enc_T_9; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_11 = has_read_req_52 ? 64'h10000000000000 : _out_read_index_enc_T_10; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_12 = has_read_req_51 ? 64'h8000000000000 : _out_read_index_enc_T_11; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_13 = has_read_req_50 ? 64'h4000000000000 : _out_read_index_enc_T_12; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_14 = has_read_req_49 ? 64'h2000000000000 : _out_read_index_enc_T_13; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_15 = has_read_req_48 ? 64'h1000000000000 : _out_read_index_enc_T_14; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_16 = has_read_req_47 ? 64'h800000000000 : _out_read_index_enc_T_15; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_17 = has_read_req_46 ? 64'h400000000000 : _out_read_index_enc_T_16; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_18 = has_read_req_45 ? 64'h200000000000 : _out_read_index_enc_T_17; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_19 = has_read_req_44 ? 64'h100000000000 : _out_read_index_enc_T_18; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_20 = has_read_req_43 ? 64'h80000000000 : _out_read_index_enc_T_19; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_21 = has_read_req_42 ? 64'h40000000000 : _out_read_index_enc_T_20; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_22 = has_read_req_41 ? 64'h20000000000 : _out_read_index_enc_T_21; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_23 = has_read_req_40 ? 64'h10000000000 : _out_read_index_enc_T_22; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_24 = has_read_req_39 ? 64'h8000000000 : _out_read_index_enc_T_23; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_25 = has_read_req_38 ? 64'h4000000000 : _out_read_index_enc_T_24; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_26 = has_read_req_37 ? 64'h2000000000 : _out_read_index_enc_T_25; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_27 = has_read_req_36 ? 64'h1000000000 : _out_read_index_enc_T_26; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_28 = has_read_req_35 ? 64'h800000000 : _out_read_index_enc_T_27; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_29 = has_read_req_34 ? 64'h400000000 : _out_read_index_enc_T_28; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_30 = has_read_req_33 ? 64'h200000000 : _out_read_index_enc_T_29; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_31 = has_read_req_32 ? 64'h100000000 : _out_read_index_enc_T_30; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_32 = has_read_req_31 ? 64'h80000000 : _out_read_index_enc_T_31; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_33 = has_read_req_30 ? 64'h40000000 : _out_read_index_enc_T_32; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_34 = has_read_req_29 ? 64'h20000000 : _out_read_index_enc_T_33; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_35 = has_read_req_28 ? 64'h10000000 : _out_read_index_enc_T_34; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_36 = has_read_req_27 ? 64'h8000000 : _out_read_index_enc_T_35; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_37 = has_read_req_26 ? 64'h4000000 : _out_read_index_enc_T_36; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_38 = has_read_req_25 ? 64'h2000000 : _out_read_index_enc_T_37; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_39 = has_read_req_24 ? 64'h1000000 : _out_read_index_enc_T_38; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_40 = has_read_req_23 ? 64'h800000 : _out_read_index_enc_T_39; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_41 = has_read_req_22 ? 64'h400000 : _out_read_index_enc_T_40; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_42 = has_read_req_21 ? 64'h200000 : _out_read_index_enc_T_41; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_43 = has_read_req_20 ? 64'h100000 : _out_read_index_enc_T_42; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_44 = has_read_req_19 ? 64'h80000 : _out_read_index_enc_T_43; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_45 = has_read_req_18 ? 64'h40000 : _out_read_index_enc_T_44; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_46 = has_read_req_17 ? 64'h20000 : _out_read_index_enc_T_45; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_47 = has_read_req_16 ? 64'h10000 : _out_read_index_enc_T_46; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_48 = has_read_req_15 ? 64'h8000 : _out_read_index_enc_T_47; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_49 = has_read_req_14 ? 64'h4000 : _out_read_index_enc_T_48; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_50 = has_read_req_13 ? 64'h2000 : _out_read_index_enc_T_49; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_51 = has_read_req_12 ? 64'h1000 : _out_read_index_enc_T_50; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_52 = has_read_req_11 ? 64'h800 : _out_read_index_enc_T_51; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_53 = has_read_req_10 ? 64'h400 : _out_read_index_enc_T_52; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_54 = has_read_req_9 ? 64'h200 : _out_read_index_enc_T_53; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_55 = has_read_req_8 ? 64'h100 : _out_read_index_enc_T_54; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_56 = has_read_req_7 ? 64'h80 : _out_read_index_enc_T_55; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_57 = has_read_req_6 ? 64'h40 : _out_read_index_enc_T_56; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_58 = has_read_req_5 ? 64'h20 : _out_read_index_enc_T_57; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_59 = has_read_req_4 ? 64'h10 : _out_read_index_enc_T_58; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_60 = has_read_req_3 ? 64'h8 : _out_read_index_enc_T_59; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_61 = has_read_req_2 ? 64'h4 : _out_read_index_enc_T_60; // @[Mux.scala 47:70]
  wire [63:0] _out_read_index_enc_T_62 = has_read_req_1 ? 64'h2 : _out_read_index_enc_T_61; // @[Mux.scala 47:70]
  wire [63:0] out_read_index_enc = has_read_req_0 ? 64'h1 : _out_read_index_enc_T_62; // @[Mux.scala 47:70]
  wire  out_read_index_0 = out_read_index_enc[0]; // @[OneHot.scala 82:30]
  wire  out_read_index_1 = out_read_index_enc[1]; // @[OneHot.scala 82:30]
  wire  out_read_index_2 = out_read_index_enc[2]; // @[OneHot.scala 82:30]
  wire  out_read_index_3 = out_read_index_enc[3]; // @[OneHot.scala 82:30]
  wire  out_read_index_4 = out_read_index_enc[4]; // @[OneHot.scala 82:30]
  wire  out_read_index_5 = out_read_index_enc[5]; // @[OneHot.scala 82:30]
  wire  out_read_index_6 = out_read_index_enc[6]; // @[OneHot.scala 82:30]
  wire  out_read_index_7 = out_read_index_enc[7]; // @[OneHot.scala 82:30]
  wire  out_read_index_8 = out_read_index_enc[8]; // @[OneHot.scala 82:30]
  wire  out_read_index_9 = out_read_index_enc[9]; // @[OneHot.scala 82:30]
  wire  out_read_index_10 = out_read_index_enc[10]; // @[OneHot.scala 82:30]
  wire  out_read_index_11 = out_read_index_enc[11]; // @[OneHot.scala 82:30]
  wire  out_read_index_12 = out_read_index_enc[12]; // @[OneHot.scala 82:30]
  wire  out_read_index_13 = out_read_index_enc[13]; // @[OneHot.scala 82:30]
  wire  out_read_index_14 = out_read_index_enc[14]; // @[OneHot.scala 82:30]
  wire  out_read_index_15 = out_read_index_enc[15]; // @[OneHot.scala 82:30]
  wire  out_read_index_16 = out_read_index_enc[16]; // @[OneHot.scala 82:30]
  wire  out_read_index_17 = out_read_index_enc[17]; // @[OneHot.scala 82:30]
  wire  out_read_index_18 = out_read_index_enc[18]; // @[OneHot.scala 82:30]
  wire  out_read_index_19 = out_read_index_enc[19]; // @[OneHot.scala 82:30]
  wire  out_read_index_20 = out_read_index_enc[20]; // @[OneHot.scala 82:30]
  wire  out_read_index_21 = out_read_index_enc[21]; // @[OneHot.scala 82:30]
  wire  out_read_index_22 = out_read_index_enc[22]; // @[OneHot.scala 82:30]
  wire  out_read_index_23 = out_read_index_enc[23]; // @[OneHot.scala 82:30]
  wire  out_read_index_24 = out_read_index_enc[24]; // @[OneHot.scala 82:30]
  wire  out_read_index_25 = out_read_index_enc[25]; // @[OneHot.scala 82:30]
  wire  out_read_index_26 = out_read_index_enc[26]; // @[OneHot.scala 82:30]
  wire  out_read_index_27 = out_read_index_enc[27]; // @[OneHot.scala 82:30]
  wire  out_read_index_28 = out_read_index_enc[28]; // @[OneHot.scala 82:30]
  wire  out_read_index_29 = out_read_index_enc[29]; // @[OneHot.scala 82:30]
  wire  out_read_index_30 = out_read_index_enc[30]; // @[OneHot.scala 82:30]
  wire  out_read_index_31 = out_read_index_enc[31]; // @[OneHot.scala 82:30]
  wire  out_read_index_32 = out_read_index_enc[32]; // @[OneHot.scala 82:30]
  wire  out_read_index_33 = out_read_index_enc[33]; // @[OneHot.scala 82:30]
  wire  out_read_index_34 = out_read_index_enc[34]; // @[OneHot.scala 82:30]
  wire  out_read_index_35 = out_read_index_enc[35]; // @[OneHot.scala 82:30]
  wire  out_read_index_36 = out_read_index_enc[36]; // @[OneHot.scala 82:30]
  wire  out_read_index_37 = out_read_index_enc[37]; // @[OneHot.scala 82:30]
  wire  out_read_index_38 = out_read_index_enc[38]; // @[OneHot.scala 82:30]
  wire  out_read_index_39 = out_read_index_enc[39]; // @[OneHot.scala 82:30]
  wire  out_read_index_40 = out_read_index_enc[40]; // @[OneHot.scala 82:30]
  wire  out_read_index_41 = out_read_index_enc[41]; // @[OneHot.scala 82:30]
  wire  out_read_index_42 = out_read_index_enc[42]; // @[OneHot.scala 82:30]
  wire  out_read_index_43 = out_read_index_enc[43]; // @[OneHot.scala 82:30]
  wire  out_read_index_44 = out_read_index_enc[44]; // @[OneHot.scala 82:30]
  wire  out_read_index_45 = out_read_index_enc[45]; // @[OneHot.scala 82:30]
  wire  out_read_index_46 = out_read_index_enc[46]; // @[OneHot.scala 82:30]
  wire  out_read_index_47 = out_read_index_enc[47]; // @[OneHot.scala 82:30]
  wire  out_read_index_48 = out_read_index_enc[48]; // @[OneHot.scala 82:30]
  wire  out_read_index_49 = out_read_index_enc[49]; // @[OneHot.scala 82:30]
  wire  out_read_index_50 = out_read_index_enc[50]; // @[OneHot.scala 82:30]
  wire  out_read_index_51 = out_read_index_enc[51]; // @[OneHot.scala 82:30]
  wire  out_read_index_52 = out_read_index_enc[52]; // @[OneHot.scala 82:30]
  wire  out_read_index_53 = out_read_index_enc[53]; // @[OneHot.scala 82:30]
  wire  out_read_index_54 = out_read_index_enc[54]; // @[OneHot.scala 82:30]
  wire  out_read_index_55 = out_read_index_enc[55]; // @[OneHot.scala 82:30]
  wire  out_read_index_56 = out_read_index_enc[56]; // @[OneHot.scala 82:30]
  wire  out_read_index_57 = out_read_index_enc[57]; // @[OneHot.scala 82:30]
  wire  out_read_index_58 = out_read_index_enc[58]; // @[OneHot.scala 82:30]
  wire  out_read_index_59 = out_read_index_enc[59]; // @[OneHot.scala 82:30]
  wire  out_read_index_60 = out_read_index_enc[60]; // @[OneHot.scala 82:30]
  wire  out_read_index_61 = out_read_index_enc[61]; // @[OneHot.scala 82:30]
  wire  out_read_index_62 = out_read_index_enc[62]; // @[OneHot.scala 82:30]
  wire  out_read_index_63 = out_read_index_enc[63]; // @[OneHot.scala 82:30]
  wire [63:0] _out_read_req_T_254 = out_read_index_0 ? mshr_0_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_255 = out_read_index_1 ? mshr_1_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_256 = out_read_index_2 ? mshr_2_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_257 = out_read_index_3 ? mshr_3_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_258 = out_read_index_4 ? mshr_4_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_259 = out_read_index_5 ? mshr_5_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_260 = out_read_index_6 ? mshr_6_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_261 = out_read_index_7 ? mshr_7_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_262 = out_read_index_8 ? mshr_8_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_263 = out_read_index_9 ? mshr_9_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_264 = out_read_index_10 ? mshr_10_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_265 = out_read_index_11 ? mshr_11_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_266 = out_read_index_12 ? mshr_12_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_267 = out_read_index_13 ? mshr_13_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_268 = out_read_index_14 ? mshr_14_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_269 = out_read_index_15 ? mshr_15_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_270 = out_read_index_16 ? mshr_16_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_271 = out_read_index_17 ? mshr_17_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_272 = out_read_index_18 ? mshr_18_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_273 = out_read_index_19 ? mshr_19_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_274 = out_read_index_20 ? mshr_20_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_275 = out_read_index_21 ? mshr_21_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_276 = out_read_index_22 ? mshr_22_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_277 = out_read_index_23 ? mshr_23_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_278 = out_read_index_24 ? mshr_24_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_279 = out_read_index_25 ? mshr_25_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_280 = out_read_index_26 ? mshr_26_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_281 = out_read_index_27 ? mshr_27_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_282 = out_read_index_28 ? mshr_28_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_283 = out_read_index_29 ? mshr_29_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_284 = out_read_index_30 ? mshr_30_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_285 = out_read_index_31 ? mshr_31_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_286 = out_read_index_32 ? mshr_32_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_287 = out_read_index_33 ? mshr_33_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_288 = out_read_index_34 ? mshr_34_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_289 = out_read_index_35 ? mshr_35_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_290 = out_read_index_36 ? mshr_36_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_291 = out_read_index_37 ? mshr_37_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_292 = out_read_index_38 ? mshr_38_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_293 = out_read_index_39 ? mshr_39_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_294 = out_read_index_40 ? mshr_40_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_295 = out_read_index_41 ? mshr_41_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_296 = out_read_index_42 ? mshr_42_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_297 = out_read_index_43 ? mshr_43_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_298 = out_read_index_44 ? mshr_44_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_299 = out_read_index_45 ? mshr_45_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_300 = out_read_index_46 ? mshr_46_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_301 = out_read_index_47 ? mshr_47_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_302 = out_read_index_48 ? mshr_48_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_303 = out_read_index_49 ? mshr_49_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_304 = out_read_index_50 ? mshr_50_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_305 = out_read_index_51 ? mshr_51_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_306 = out_read_index_52 ? mshr_52_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_307 = out_read_index_53 ? mshr_53_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_308 = out_read_index_54 ? mshr_54_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_309 = out_read_index_55 ? mshr_55_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_310 = out_read_index_56 ? mshr_56_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_311 = out_read_index_57 ? mshr_57_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_312 = out_read_index_58 ? mshr_58_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_313 = out_read_index_59 ? mshr_59_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_314 = out_read_index_60 ? mshr_60_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_315 = out_read_index_61 ? mshr_61_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_316 = out_read_index_62 ? mshr_62_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_317 = out_read_index_63 ? mshr_63_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_318 = _out_read_req_T_254 | _out_read_req_T_255; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_319 = _out_read_req_T_318 | _out_read_req_T_256; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_320 = _out_read_req_T_319 | _out_read_req_T_257; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_321 = _out_read_req_T_320 | _out_read_req_T_258; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_322 = _out_read_req_T_321 | _out_read_req_T_259; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_323 = _out_read_req_T_322 | _out_read_req_T_260; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_324 = _out_read_req_T_323 | _out_read_req_T_261; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_325 = _out_read_req_T_324 | _out_read_req_T_262; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_326 = _out_read_req_T_325 | _out_read_req_T_263; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_327 = _out_read_req_T_326 | _out_read_req_T_264; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_328 = _out_read_req_T_327 | _out_read_req_T_265; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_329 = _out_read_req_T_328 | _out_read_req_T_266; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_330 = _out_read_req_T_329 | _out_read_req_T_267; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_331 = _out_read_req_T_330 | _out_read_req_T_268; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_332 = _out_read_req_T_331 | _out_read_req_T_269; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_333 = _out_read_req_T_332 | _out_read_req_T_270; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_334 = _out_read_req_T_333 | _out_read_req_T_271; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_335 = _out_read_req_T_334 | _out_read_req_T_272; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_336 = _out_read_req_T_335 | _out_read_req_T_273; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_337 = _out_read_req_T_336 | _out_read_req_T_274; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_338 = _out_read_req_T_337 | _out_read_req_T_275; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_339 = _out_read_req_T_338 | _out_read_req_T_276; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_340 = _out_read_req_T_339 | _out_read_req_T_277; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_341 = _out_read_req_T_340 | _out_read_req_T_278; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_342 = _out_read_req_T_341 | _out_read_req_T_279; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_343 = _out_read_req_T_342 | _out_read_req_T_280; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_344 = _out_read_req_T_343 | _out_read_req_T_281; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_345 = _out_read_req_T_344 | _out_read_req_T_282; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_346 = _out_read_req_T_345 | _out_read_req_T_283; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_347 = _out_read_req_T_346 | _out_read_req_T_284; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_348 = _out_read_req_T_347 | _out_read_req_T_285; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_349 = _out_read_req_T_348 | _out_read_req_T_286; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_350 = _out_read_req_T_349 | _out_read_req_T_287; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_351 = _out_read_req_T_350 | _out_read_req_T_288; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_352 = _out_read_req_T_351 | _out_read_req_T_289; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_353 = _out_read_req_T_352 | _out_read_req_T_290; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_354 = _out_read_req_T_353 | _out_read_req_T_291; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_355 = _out_read_req_T_354 | _out_read_req_T_292; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_356 = _out_read_req_T_355 | _out_read_req_T_293; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_357 = _out_read_req_T_356 | _out_read_req_T_294; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_358 = _out_read_req_T_357 | _out_read_req_T_295; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_359 = _out_read_req_T_358 | _out_read_req_T_296; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_360 = _out_read_req_T_359 | _out_read_req_T_297; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_361 = _out_read_req_T_360 | _out_read_req_T_298; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_362 = _out_read_req_T_361 | _out_read_req_T_299; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_363 = _out_read_req_T_362 | _out_read_req_T_300; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_364 = _out_read_req_T_363 | _out_read_req_T_301; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_365 = _out_read_req_T_364 | _out_read_req_T_302; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_366 = _out_read_req_T_365 | _out_read_req_T_303; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_367 = _out_read_req_T_366 | _out_read_req_T_304; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_368 = _out_read_req_T_367 | _out_read_req_T_305; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_369 = _out_read_req_T_368 | _out_read_req_T_306; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_370 = _out_read_req_T_369 | _out_read_req_T_307; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_371 = _out_read_req_T_370 | _out_read_req_T_308; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_372 = _out_read_req_T_371 | _out_read_req_T_309; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_373 = _out_read_req_T_372 | _out_read_req_T_310; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_374 = _out_read_req_T_373 | _out_read_req_T_311; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_375 = _out_read_req_T_374 | _out_read_req_T_312; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_376 = _out_read_req_T_375 | _out_read_req_T_313; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_377 = _out_read_req_T_376 | _out_read_req_T_314; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_378 = _out_read_req_T_377 | _out_read_req_T_315; // @[Mux.scala 27:73]
  wire [63:0] _out_read_req_T_379 = _out_read_req_T_378 | _out_read_req_T_316; // @[Mux.scala 27:73]
  wire [63:0] out_read_req_addr = _out_read_req_T_379 | _out_read_req_T_317; // @[Mux.scala 27:73]
  wire [7:0] bundleOut_0_arvalid_lo_lo_lo = {has_read_req_7,has_read_req_6,has_read_req_5,has_read_req_4,has_read_req_3
    ,has_read_req_2,has_read_req_1,has_read_req_0}; // @[AXI4FakeDMA.scala 187:34]
  wire [15:0] bundleOut_0_arvalid_lo_lo = {has_read_req_15,has_read_req_14,has_read_req_13,has_read_req_12,
    has_read_req_11,has_read_req_10,has_read_req_9,has_read_req_8,bundleOut_0_arvalid_lo_lo_lo}; // @[AXI4FakeDMA.scala 187:34]
  wire [7:0] bundleOut_0_arvalid_lo_hi_lo = {has_read_req_23,has_read_req_22,has_read_req_21,has_read_req_20,
    has_read_req_19,has_read_req_18,has_read_req_17,has_read_req_16}; // @[AXI4FakeDMA.scala 187:34]
  wire [31:0] bundleOut_0_arvalid_lo = {has_read_req_31,has_read_req_30,has_read_req_29,has_read_req_28,has_read_req_27
    ,has_read_req_26,has_read_req_25,has_read_req_24,bundleOut_0_arvalid_lo_hi_lo,bundleOut_0_arvalid_lo_lo}; // @[AXI4FakeDMA.scala 187:34]
  wire [7:0] bundleOut_0_arvalid_hi_lo_lo = {has_read_req_39,has_read_req_38,has_read_req_37,has_read_req_36,
    has_read_req_35,has_read_req_34,has_read_req_33,has_read_req_32}; // @[AXI4FakeDMA.scala 187:34]
  wire [15:0] bundleOut_0_arvalid_hi_lo = {has_read_req_47,has_read_req_46,has_read_req_45,has_read_req_44,
    has_read_req_43,has_read_req_42,has_read_req_41,has_read_req_40,bundleOut_0_arvalid_hi_lo_lo}; // @[AXI4FakeDMA.scala 187:34]
  wire [7:0] bundleOut_0_arvalid_hi_hi_lo = {has_read_req_55,has_read_req_54,has_read_req_53,has_read_req_52,
    has_read_req_51,has_read_req_50,has_read_req_49,has_read_req_48}; // @[AXI4FakeDMA.scala 187:34]
  wire [31:0] bundleOut_0_arvalid_hi = {has_read_req_63,has_read_req_62,has_read_req_61,has_read_req_60,has_read_req_59
    ,has_read_req_58,has_read_req_57,has_read_req_56,bundleOut_0_arvalid_hi_hi_lo,bundleOut_0_arvalid_hi_lo}; // @[AXI4FakeDMA.scala 187:34]
  wire [63:0] _bundleOut_0_arvalid_T = {bundleOut_0_arvalid_hi,bundleOut_0_arvalid_lo}; // @[AXI4FakeDMA.scala 187:34]
  wire  out_arvalid = |_bundleOut_0_arvalid_T; // @[AXI4FakeDMA.scala 187:41]
  wire [7:0] bundleOut_0_arid_lo_lo_lo = {out_read_index_7,out_read_index_6,out_read_index_5,out_read_index_4,
    out_read_index_3,out_read_index_2,out_read_index_1,out_read_index_0}; // @[Cat.scala 31:58]
  wire [15:0] bundleOut_0_arid_lo_lo = {out_read_index_15,out_read_index_14,out_read_index_13,out_read_index_12,
    out_read_index_11,out_read_index_10,out_read_index_9,out_read_index_8,bundleOut_0_arid_lo_lo_lo}; // @[Cat.scala 31:58]
  wire [7:0] bundleOut_0_arid_lo_hi_lo = {out_read_index_23,out_read_index_22,out_read_index_21,out_read_index_20,
    out_read_index_19,out_read_index_18,out_read_index_17,out_read_index_16}; // @[Cat.scala 31:58]
  wire [31:0] bundleOut_0_arid_lo = {out_read_index_31,out_read_index_30,out_read_index_29,out_read_index_28,
    out_read_index_27,out_read_index_26,out_read_index_25,out_read_index_24,bundleOut_0_arid_lo_hi_lo,
    bundleOut_0_arid_lo_lo}; // @[Cat.scala 31:58]
  wire [7:0] bundleOut_0_arid_hi_lo_lo = {out_read_index_39,out_read_index_38,out_read_index_37,out_read_index_36,
    out_read_index_35,out_read_index_34,out_read_index_33,out_read_index_32}; // @[Cat.scala 31:58]
  wire [15:0] bundleOut_0_arid_hi_lo = {out_read_index_47,out_read_index_46,out_read_index_45,out_read_index_44,
    out_read_index_43,out_read_index_42,out_read_index_41,out_read_index_40,bundleOut_0_arid_hi_lo_lo}; // @[Cat.scala 31:58]
  wire [7:0] bundleOut_0_arid_hi_hi_lo = {out_read_index_55,out_read_index_54,out_read_index_53,out_read_index_52,
    out_read_index_51,out_read_index_50,out_read_index_49,out_read_index_48}; // @[Cat.scala 31:58]
  wire [31:0] bundleOut_0_arid_hi = {out_read_index_63,out_read_index_62,out_read_index_61,out_read_index_60,
    out_read_index_59,out_read_index_58,out_read_index_57,out_read_index_56,bundleOut_0_arid_hi_hi_lo,
    bundleOut_0_arid_hi_lo}; // @[Cat.scala 31:58]
  wire [63:0] _bundleOut_0_arid_T = {bundleOut_0_arid_hi,bundleOut_0_arid_lo}; // @[Cat.scala 31:58]
  wire [31:0] bundleOut_0_arid_hi_1 = _bundleOut_0_arid_T[63:32]; // @[OneHot.scala 30:18]
  wire [31:0] bundleOut_0_arid_lo_1 = _bundleOut_0_arid_T[31:0]; // @[OneHot.scala 31:18]
  wire  _bundleOut_0_arid_T_1 = |bundleOut_0_arid_hi_1; // @[OneHot.scala 32:14]
  wire [31:0] _bundleOut_0_arid_T_2 = bundleOut_0_arid_hi_1 | bundleOut_0_arid_lo_1; // @[OneHot.scala 32:28]
  wire [15:0] bundleOut_0_arid_hi_2 = _bundleOut_0_arid_T_2[31:16]; // @[OneHot.scala 30:18]
  wire [15:0] bundleOut_0_arid_lo_2 = _bundleOut_0_arid_T_2[15:0]; // @[OneHot.scala 31:18]
  wire  _bundleOut_0_arid_T_3 = |bundleOut_0_arid_hi_2; // @[OneHot.scala 32:14]
  wire [15:0] _bundleOut_0_arid_T_4 = bundleOut_0_arid_hi_2 | bundleOut_0_arid_lo_2; // @[OneHot.scala 32:28]
  wire [7:0] bundleOut_0_arid_hi_3 = _bundleOut_0_arid_T_4[15:8]; // @[OneHot.scala 30:18]
  wire [7:0] bundleOut_0_arid_lo_3 = _bundleOut_0_arid_T_4[7:0]; // @[OneHot.scala 31:18]
  wire  _bundleOut_0_arid_T_5 = |bundleOut_0_arid_hi_3; // @[OneHot.scala 32:14]
  wire [7:0] _bundleOut_0_arid_T_6 = bundleOut_0_arid_hi_3 | bundleOut_0_arid_lo_3; // @[OneHot.scala 32:28]
  wire [3:0] bundleOut_0_arid_hi_4 = _bundleOut_0_arid_T_6[7:4]; // @[OneHot.scala 30:18]
  wire [3:0] bundleOut_0_arid_lo_4 = _bundleOut_0_arid_T_6[3:0]; // @[OneHot.scala 31:18]
  wire  _bundleOut_0_arid_T_7 = |bundleOut_0_arid_hi_4; // @[OneHot.scala 32:14]
  wire [3:0] _bundleOut_0_arid_T_8 = bundleOut_0_arid_hi_4 | bundleOut_0_arid_lo_4; // @[OneHot.scala 32:28]
  wire [1:0] bundleOut_0_arid_hi_5 = _bundleOut_0_arid_T_8[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] bundleOut_0_arid_lo_5 = _bundleOut_0_arid_T_8[1:0]; // @[OneHot.scala 31:18]
  wire  _bundleOut_0_arid_T_9 = |bundleOut_0_arid_hi_5; // @[OneHot.scala 32:14]
  wire [1:0] _bundleOut_0_arid_T_10 = bundleOut_0_arid_hi_5 | bundleOut_0_arid_lo_5; // @[OneHot.scala 32:28]
  wire [5:0] _bundleOut_0_arid_T_16 = {_bundleOut_0_arid_T_1,_bundleOut_0_arid_T_3,
    _bundleOut_0_arid_T_5,_bundleOut_0_arid_T_7,_bundleOut_0_arid_T_9,_bundleOut_0_arid_T_10[1]}
    ; // @[Cat.scala 31:58]
  wire  has_write_req_0 = mshr_0_io_master_req_valid & mshr_0_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_1 = mshr_1_io_master_req_valid & mshr_1_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_2 = mshr_2_io_master_req_valid & mshr_2_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_3 = mshr_3_io_master_req_valid & mshr_3_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_4 = mshr_4_io_master_req_valid & mshr_4_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_5 = mshr_5_io_master_req_valid & mshr_5_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_6 = mshr_6_io_master_req_valid & mshr_6_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_7 = mshr_7_io_master_req_valid & mshr_7_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_8 = mshr_8_io_master_req_valid & mshr_8_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_9 = mshr_9_io_master_req_valid & mshr_9_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_10 = mshr_10_io_master_req_valid & mshr_10_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_11 = mshr_11_io_master_req_valid & mshr_11_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_12 = mshr_12_io_master_req_valid & mshr_12_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_13 = mshr_13_io_master_req_valid & mshr_13_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_14 = mshr_14_io_master_req_valid & mshr_14_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_15 = mshr_15_io_master_req_valid & mshr_15_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_16 = mshr_16_io_master_req_valid & mshr_16_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_17 = mshr_17_io_master_req_valid & mshr_17_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_18 = mshr_18_io_master_req_valid & mshr_18_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_19 = mshr_19_io_master_req_valid & mshr_19_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_20 = mshr_20_io_master_req_valid & mshr_20_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_21 = mshr_21_io_master_req_valid & mshr_21_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_22 = mshr_22_io_master_req_valid & mshr_22_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_23 = mshr_23_io_master_req_valid & mshr_23_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_24 = mshr_24_io_master_req_valid & mshr_24_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_25 = mshr_25_io_master_req_valid & mshr_25_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_26 = mshr_26_io_master_req_valid & mshr_26_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_27 = mshr_27_io_master_req_valid & mshr_27_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_28 = mshr_28_io_master_req_valid & mshr_28_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_29 = mshr_29_io_master_req_valid & mshr_29_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_30 = mshr_30_io_master_req_valid & mshr_30_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_31 = mshr_31_io_master_req_valid & mshr_31_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_32 = mshr_32_io_master_req_valid & mshr_32_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_33 = mshr_33_io_master_req_valid & mshr_33_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_34 = mshr_34_io_master_req_valid & mshr_34_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_35 = mshr_35_io_master_req_valid & mshr_35_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_36 = mshr_36_io_master_req_valid & mshr_36_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_37 = mshr_37_io_master_req_valid & mshr_37_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_38 = mshr_38_io_master_req_valid & mshr_38_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_39 = mshr_39_io_master_req_valid & mshr_39_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_40 = mshr_40_io_master_req_valid & mshr_40_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_41 = mshr_41_io_master_req_valid & mshr_41_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_42 = mshr_42_io_master_req_valid & mshr_42_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_43 = mshr_43_io_master_req_valid & mshr_43_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_44 = mshr_44_io_master_req_valid & mshr_44_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_45 = mshr_45_io_master_req_valid & mshr_45_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_46 = mshr_46_io_master_req_valid & mshr_46_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_47 = mshr_47_io_master_req_valid & mshr_47_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_48 = mshr_48_io_master_req_valid & mshr_48_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_49 = mshr_49_io_master_req_valid & mshr_49_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_50 = mshr_50_io_master_req_valid & mshr_50_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_51 = mshr_51_io_master_req_valid & mshr_51_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_52 = mshr_52_io_master_req_valid & mshr_52_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_53 = mshr_53_io_master_req_valid & mshr_53_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_54 = mshr_54_io_master_req_valid & mshr_54_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_55 = mshr_55_io_master_req_valid & mshr_55_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_56 = mshr_56_io_master_req_valid & mshr_56_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_57 = mshr_57_io_master_req_valid & mshr_57_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_58 = mshr_58_io_master_req_valid & mshr_58_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_59 = mshr_59_io_master_req_valid & mshr_59_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_60 = mshr_60_io_master_req_valid & mshr_60_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_61 = mshr_61_io_master_req_valid & mshr_61_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_62 = mshr_62_io_master_req_valid & mshr_62_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire  has_write_req_63 = mshr_63_io_master_req_valid & mshr_63_io_master_req_is_write; // @[AXI4FakeDMA.scala 132:49]
  wire [63:0] _out_write_index_enc_T = has_write_req_63 ? 64'h8000000000000000 : 64'h0; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_1 = has_write_req_62 ? 64'h4000000000000000 : _out_write_index_enc_T; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_2 = has_write_req_61 ? 64'h2000000000000000 : _out_write_index_enc_T_1; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_3 = has_write_req_60 ? 64'h1000000000000000 : _out_write_index_enc_T_2; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_4 = has_write_req_59 ? 64'h800000000000000 : _out_write_index_enc_T_3; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_5 = has_write_req_58 ? 64'h400000000000000 : _out_write_index_enc_T_4; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_6 = has_write_req_57 ? 64'h200000000000000 : _out_write_index_enc_T_5; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_7 = has_write_req_56 ? 64'h100000000000000 : _out_write_index_enc_T_6; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_8 = has_write_req_55 ? 64'h80000000000000 : _out_write_index_enc_T_7; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_9 = has_write_req_54 ? 64'h40000000000000 : _out_write_index_enc_T_8; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_10 = has_write_req_53 ? 64'h20000000000000 : _out_write_index_enc_T_9; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_11 = has_write_req_52 ? 64'h10000000000000 : _out_write_index_enc_T_10; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_12 = has_write_req_51 ? 64'h8000000000000 : _out_write_index_enc_T_11; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_13 = has_write_req_50 ? 64'h4000000000000 : _out_write_index_enc_T_12; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_14 = has_write_req_49 ? 64'h2000000000000 : _out_write_index_enc_T_13; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_15 = has_write_req_48 ? 64'h1000000000000 : _out_write_index_enc_T_14; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_16 = has_write_req_47 ? 64'h800000000000 : _out_write_index_enc_T_15; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_17 = has_write_req_46 ? 64'h400000000000 : _out_write_index_enc_T_16; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_18 = has_write_req_45 ? 64'h200000000000 : _out_write_index_enc_T_17; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_19 = has_write_req_44 ? 64'h100000000000 : _out_write_index_enc_T_18; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_20 = has_write_req_43 ? 64'h80000000000 : _out_write_index_enc_T_19; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_21 = has_write_req_42 ? 64'h40000000000 : _out_write_index_enc_T_20; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_22 = has_write_req_41 ? 64'h20000000000 : _out_write_index_enc_T_21; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_23 = has_write_req_40 ? 64'h10000000000 : _out_write_index_enc_T_22; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_24 = has_write_req_39 ? 64'h8000000000 : _out_write_index_enc_T_23; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_25 = has_write_req_38 ? 64'h4000000000 : _out_write_index_enc_T_24; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_26 = has_write_req_37 ? 64'h2000000000 : _out_write_index_enc_T_25; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_27 = has_write_req_36 ? 64'h1000000000 : _out_write_index_enc_T_26; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_28 = has_write_req_35 ? 64'h800000000 : _out_write_index_enc_T_27; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_29 = has_write_req_34 ? 64'h400000000 : _out_write_index_enc_T_28; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_30 = has_write_req_33 ? 64'h200000000 : _out_write_index_enc_T_29; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_31 = has_write_req_32 ? 64'h100000000 : _out_write_index_enc_T_30; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_32 = has_write_req_31 ? 64'h80000000 : _out_write_index_enc_T_31; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_33 = has_write_req_30 ? 64'h40000000 : _out_write_index_enc_T_32; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_34 = has_write_req_29 ? 64'h20000000 : _out_write_index_enc_T_33; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_35 = has_write_req_28 ? 64'h10000000 : _out_write_index_enc_T_34; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_36 = has_write_req_27 ? 64'h8000000 : _out_write_index_enc_T_35; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_37 = has_write_req_26 ? 64'h4000000 : _out_write_index_enc_T_36; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_38 = has_write_req_25 ? 64'h2000000 : _out_write_index_enc_T_37; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_39 = has_write_req_24 ? 64'h1000000 : _out_write_index_enc_T_38; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_40 = has_write_req_23 ? 64'h800000 : _out_write_index_enc_T_39; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_41 = has_write_req_22 ? 64'h400000 : _out_write_index_enc_T_40; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_42 = has_write_req_21 ? 64'h200000 : _out_write_index_enc_T_41; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_43 = has_write_req_20 ? 64'h100000 : _out_write_index_enc_T_42; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_44 = has_write_req_19 ? 64'h80000 : _out_write_index_enc_T_43; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_45 = has_write_req_18 ? 64'h40000 : _out_write_index_enc_T_44; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_46 = has_write_req_17 ? 64'h20000 : _out_write_index_enc_T_45; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_47 = has_write_req_16 ? 64'h10000 : _out_write_index_enc_T_46; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_48 = has_write_req_15 ? 64'h8000 : _out_write_index_enc_T_47; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_49 = has_write_req_14 ? 64'h4000 : _out_write_index_enc_T_48; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_50 = has_write_req_13 ? 64'h2000 : _out_write_index_enc_T_49; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_51 = has_write_req_12 ? 64'h1000 : _out_write_index_enc_T_50; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_52 = has_write_req_11 ? 64'h800 : _out_write_index_enc_T_51; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_53 = has_write_req_10 ? 64'h400 : _out_write_index_enc_T_52; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_54 = has_write_req_9 ? 64'h200 : _out_write_index_enc_T_53; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_55 = has_write_req_8 ? 64'h100 : _out_write_index_enc_T_54; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_56 = has_write_req_7 ? 64'h80 : _out_write_index_enc_T_55; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_57 = has_write_req_6 ? 64'h40 : _out_write_index_enc_T_56; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_58 = has_write_req_5 ? 64'h20 : _out_write_index_enc_T_57; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_59 = has_write_req_4 ? 64'h10 : _out_write_index_enc_T_58; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_60 = has_write_req_3 ? 64'h8 : _out_write_index_enc_T_59; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_61 = has_write_req_2 ? 64'h4 : _out_write_index_enc_T_60; // @[Mux.scala 47:70]
  wire [63:0] _out_write_index_enc_T_62 = has_write_req_1 ? 64'h2 : _out_write_index_enc_T_61; // @[Mux.scala 47:70]
  wire [63:0] out_write_index_enc = has_write_req_0 ? 64'h1 : _out_write_index_enc_T_62; // @[Mux.scala 47:70]
  wire  out_write_index_0 = out_write_index_enc[0]; // @[OneHot.scala 82:30]
  wire  out_write_index_1 = out_write_index_enc[1]; // @[OneHot.scala 82:30]
  wire  out_write_index_2 = out_write_index_enc[2]; // @[OneHot.scala 82:30]
  wire  out_write_index_3 = out_write_index_enc[3]; // @[OneHot.scala 82:30]
  wire  out_write_index_4 = out_write_index_enc[4]; // @[OneHot.scala 82:30]
  wire  out_write_index_5 = out_write_index_enc[5]; // @[OneHot.scala 82:30]
  wire  out_write_index_6 = out_write_index_enc[6]; // @[OneHot.scala 82:30]
  wire  out_write_index_7 = out_write_index_enc[7]; // @[OneHot.scala 82:30]
  wire  out_write_index_8 = out_write_index_enc[8]; // @[OneHot.scala 82:30]
  wire  out_write_index_9 = out_write_index_enc[9]; // @[OneHot.scala 82:30]
  wire  out_write_index_10 = out_write_index_enc[10]; // @[OneHot.scala 82:30]
  wire  out_write_index_11 = out_write_index_enc[11]; // @[OneHot.scala 82:30]
  wire  out_write_index_12 = out_write_index_enc[12]; // @[OneHot.scala 82:30]
  wire  out_write_index_13 = out_write_index_enc[13]; // @[OneHot.scala 82:30]
  wire  out_write_index_14 = out_write_index_enc[14]; // @[OneHot.scala 82:30]
  wire  out_write_index_15 = out_write_index_enc[15]; // @[OneHot.scala 82:30]
  wire  out_write_index_16 = out_write_index_enc[16]; // @[OneHot.scala 82:30]
  wire  out_write_index_17 = out_write_index_enc[17]; // @[OneHot.scala 82:30]
  wire  out_write_index_18 = out_write_index_enc[18]; // @[OneHot.scala 82:30]
  wire  out_write_index_19 = out_write_index_enc[19]; // @[OneHot.scala 82:30]
  wire  out_write_index_20 = out_write_index_enc[20]; // @[OneHot.scala 82:30]
  wire  out_write_index_21 = out_write_index_enc[21]; // @[OneHot.scala 82:30]
  wire  out_write_index_22 = out_write_index_enc[22]; // @[OneHot.scala 82:30]
  wire  out_write_index_23 = out_write_index_enc[23]; // @[OneHot.scala 82:30]
  wire  out_write_index_24 = out_write_index_enc[24]; // @[OneHot.scala 82:30]
  wire  out_write_index_25 = out_write_index_enc[25]; // @[OneHot.scala 82:30]
  wire  out_write_index_26 = out_write_index_enc[26]; // @[OneHot.scala 82:30]
  wire  out_write_index_27 = out_write_index_enc[27]; // @[OneHot.scala 82:30]
  wire  out_write_index_28 = out_write_index_enc[28]; // @[OneHot.scala 82:30]
  wire  out_write_index_29 = out_write_index_enc[29]; // @[OneHot.scala 82:30]
  wire  out_write_index_30 = out_write_index_enc[30]; // @[OneHot.scala 82:30]
  wire  out_write_index_31 = out_write_index_enc[31]; // @[OneHot.scala 82:30]
  wire  out_write_index_32 = out_write_index_enc[32]; // @[OneHot.scala 82:30]
  wire  out_write_index_33 = out_write_index_enc[33]; // @[OneHot.scala 82:30]
  wire  out_write_index_34 = out_write_index_enc[34]; // @[OneHot.scala 82:30]
  wire  out_write_index_35 = out_write_index_enc[35]; // @[OneHot.scala 82:30]
  wire  out_write_index_36 = out_write_index_enc[36]; // @[OneHot.scala 82:30]
  wire  out_write_index_37 = out_write_index_enc[37]; // @[OneHot.scala 82:30]
  wire  out_write_index_38 = out_write_index_enc[38]; // @[OneHot.scala 82:30]
  wire  out_write_index_39 = out_write_index_enc[39]; // @[OneHot.scala 82:30]
  wire  out_write_index_40 = out_write_index_enc[40]; // @[OneHot.scala 82:30]
  wire  out_write_index_41 = out_write_index_enc[41]; // @[OneHot.scala 82:30]
  wire  out_write_index_42 = out_write_index_enc[42]; // @[OneHot.scala 82:30]
  wire  out_write_index_43 = out_write_index_enc[43]; // @[OneHot.scala 82:30]
  wire  out_write_index_44 = out_write_index_enc[44]; // @[OneHot.scala 82:30]
  wire  out_write_index_45 = out_write_index_enc[45]; // @[OneHot.scala 82:30]
  wire  out_write_index_46 = out_write_index_enc[46]; // @[OneHot.scala 82:30]
  wire  out_write_index_47 = out_write_index_enc[47]; // @[OneHot.scala 82:30]
  wire  out_write_index_48 = out_write_index_enc[48]; // @[OneHot.scala 82:30]
  wire  out_write_index_49 = out_write_index_enc[49]; // @[OneHot.scala 82:30]
  wire  out_write_index_50 = out_write_index_enc[50]; // @[OneHot.scala 82:30]
  wire  out_write_index_51 = out_write_index_enc[51]; // @[OneHot.scala 82:30]
  wire  out_write_index_52 = out_write_index_enc[52]; // @[OneHot.scala 82:30]
  wire  out_write_index_53 = out_write_index_enc[53]; // @[OneHot.scala 82:30]
  wire  out_write_index_54 = out_write_index_enc[54]; // @[OneHot.scala 82:30]
  wire  out_write_index_55 = out_write_index_enc[55]; // @[OneHot.scala 82:30]
  wire  out_write_index_56 = out_write_index_enc[56]; // @[OneHot.scala 82:30]
  wire  out_write_index_57 = out_write_index_enc[57]; // @[OneHot.scala 82:30]
  wire  out_write_index_58 = out_write_index_enc[58]; // @[OneHot.scala 82:30]
  wire  out_write_index_59 = out_write_index_enc[59]; // @[OneHot.scala 82:30]
  wire  out_write_index_60 = out_write_index_enc[60]; // @[OneHot.scala 82:30]
  wire  out_write_index_61 = out_write_index_enc[61]; // @[OneHot.scala 82:30]
  wire  out_write_index_62 = out_write_index_enc[62]; // @[OneHot.scala 82:30]
  wire  out_write_index_63 = out_write_index_enc[63]; // @[OneHot.scala 82:30]
  wire [511:0] _out_write_req_T = out_write_index_0 ? mshr_0_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_1 = out_write_index_1 ? mshr_1_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_2 = out_write_index_2 ? mshr_2_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_3 = out_write_index_3 ? mshr_3_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_4 = out_write_index_4 ? mshr_4_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_5 = out_write_index_5 ? mshr_5_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_6 = out_write_index_6 ? mshr_6_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_7 = out_write_index_7 ? mshr_7_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_8 = out_write_index_8 ? mshr_8_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_9 = out_write_index_9 ? mshr_9_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_10 = out_write_index_10 ? mshr_10_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_11 = out_write_index_11 ? mshr_11_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_12 = out_write_index_12 ? mshr_12_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_13 = out_write_index_13 ? mshr_13_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_14 = out_write_index_14 ? mshr_14_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_15 = out_write_index_15 ? mshr_15_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_16 = out_write_index_16 ? mshr_16_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_17 = out_write_index_17 ? mshr_17_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_18 = out_write_index_18 ? mshr_18_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_19 = out_write_index_19 ? mshr_19_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_20 = out_write_index_20 ? mshr_20_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_21 = out_write_index_21 ? mshr_21_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_22 = out_write_index_22 ? mshr_22_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_23 = out_write_index_23 ? mshr_23_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_24 = out_write_index_24 ? mshr_24_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_25 = out_write_index_25 ? mshr_25_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_26 = out_write_index_26 ? mshr_26_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_27 = out_write_index_27 ? mshr_27_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_28 = out_write_index_28 ? mshr_28_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_29 = out_write_index_29 ? mshr_29_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_30 = out_write_index_30 ? mshr_30_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_31 = out_write_index_31 ? mshr_31_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_32 = out_write_index_32 ? mshr_32_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_33 = out_write_index_33 ? mshr_33_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_34 = out_write_index_34 ? mshr_34_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_35 = out_write_index_35 ? mshr_35_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_36 = out_write_index_36 ? mshr_36_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_37 = out_write_index_37 ? mshr_37_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_38 = out_write_index_38 ? mshr_38_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_39 = out_write_index_39 ? mshr_39_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_40 = out_write_index_40 ? mshr_40_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_41 = out_write_index_41 ? mshr_41_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_42 = out_write_index_42 ? mshr_42_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_43 = out_write_index_43 ? mshr_43_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_44 = out_write_index_44 ? mshr_44_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_45 = out_write_index_45 ? mshr_45_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_46 = out_write_index_46 ? mshr_46_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_47 = out_write_index_47 ? mshr_47_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_48 = out_write_index_48 ? mshr_48_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_49 = out_write_index_49 ? mshr_49_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_50 = out_write_index_50 ? mshr_50_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_51 = out_write_index_51 ? mshr_51_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_52 = out_write_index_52 ? mshr_52_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_53 = out_write_index_53 ? mshr_53_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_54 = out_write_index_54 ? mshr_54_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_55 = out_write_index_55 ? mshr_55_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_56 = out_write_index_56 ? mshr_56_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_57 = out_write_index_57 ? mshr_57_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_58 = out_write_index_58 ? mshr_58_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_59 = out_write_index_59 ? mshr_59_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_60 = out_write_index_60 ? mshr_60_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_61 = out_write_index_61 ? mshr_61_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_62 = out_write_index_62 ? mshr_62_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_63 = out_write_index_63 ? mshr_63_io_master_req_data : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_64 = _out_write_req_T | _out_write_req_T_1; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_65 = _out_write_req_T_64 | _out_write_req_T_2; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_66 = _out_write_req_T_65 | _out_write_req_T_3; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_67 = _out_write_req_T_66 | _out_write_req_T_4; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_68 = _out_write_req_T_67 | _out_write_req_T_5; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_69 = _out_write_req_T_68 | _out_write_req_T_6; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_70 = _out_write_req_T_69 | _out_write_req_T_7; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_71 = _out_write_req_T_70 | _out_write_req_T_8; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_72 = _out_write_req_T_71 | _out_write_req_T_9; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_73 = _out_write_req_T_72 | _out_write_req_T_10; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_74 = _out_write_req_T_73 | _out_write_req_T_11; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_75 = _out_write_req_T_74 | _out_write_req_T_12; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_76 = _out_write_req_T_75 | _out_write_req_T_13; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_77 = _out_write_req_T_76 | _out_write_req_T_14; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_78 = _out_write_req_T_77 | _out_write_req_T_15; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_79 = _out_write_req_T_78 | _out_write_req_T_16; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_80 = _out_write_req_T_79 | _out_write_req_T_17; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_81 = _out_write_req_T_80 | _out_write_req_T_18; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_82 = _out_write_req_T_81 | _out_write_req_T_19; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_83 = _out_write_req_T_82 | _out_write_req_T_20; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_84 = _out_write_req_T_83 | _out_write_req_T_21; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_85 = _out_write_req_T_84 | _out_write_req_T_22; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_86 = _out_write_req_T_85 | _out_write_req_T_23; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_87 = _out_write_req_T_86 | _out_write_req_T_24; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_88 = _out_write_req_T_87 | _out_write_req_T_25; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_89 = _out_write_req_T_88 | _out_write_req_T_26; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_90 = _out_write_req_T_89 | _out_write_req_T_27; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_91 = _out_write_req_T_90 | _out_write_req_T_28; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_92 = _out_write_req_T_91 | _out_write_req_T_29; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_93 = _out_write_req_T_92 | _out_write_req_T_30; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_94 = _out_write_req_T_93 | _out_write_req_T_31; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_95 = _out_write_req_T_94 | _out_write_req_T_32; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_96 = _out_write_req_T_95 | _out_write_req_T_33; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_97 = _out_write_req_T_96 | _out_write_req_T_34; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_98 = _out_write_req_T_97 | _out_write_req_T_35; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_99 = _out_write_req_T_98 | _out_write_req_T_36; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_100 = _out_write_req_T_99 | _out_write_req_T_37; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_101 = _out_write_req_T_100 | _out_write_req_T_38; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_102 = _out_write_req_T_101 | _out_write_req_T_39; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_103 = _out_write_req_T_102 | _out_write_req_T_40; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_104 = _out_write_req_T_103 | _out_write_req_T_41; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_105 = _out_write_req_T_104 | _out_write_req_T_42; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_106 = _out_write_req_T_105 | _out_write_req_T_43; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_107 = _out_write_req_T_106 | _out_write_req_T_44; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_108 = _out_write_req_T_107 | _out_write_req_T_45; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_109 = _out_write_req_T_108 | _out_write_req_T_46; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_110 = _out_write_req_T_109 | _out_write_req_T_47; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_111 = _out_write_req_T_110 | _out_write_req_T_48; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_112 = _out_write_req_T_111 | _out_write_req_T_49; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_113 = _out_write_req_T_112 | _out_write_req_T_50; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_114 = _out_write_req_T_113 | _out_write_req_T_51; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_115 = _out_write_req_T_114 | _out_write_req_T_52; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_116 = _out_write_req_T_115 | _out_write_req_T_53; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_117 = _out_write_req_T_116 | _out_write_req_T_54; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_118 = _out_write_req_T_117 | _out_write_req_T_55; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_119 = _out_write_req_T_118 | _out_write_req_T_56; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_120 = _out_write_req_T_119 | _out_write_req_T_57; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_121 = _out_write_req_T_120 | _out_write_req_T_58; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_122 = _out_write_req_T_121 | _out_write_req_T_59; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_123 = _out_write_req_T_122 | _out_write_req_T_60; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_124 = _out_write_req_T_123 | _out_write_req_T_61; // @[Mux.scala 27:73]
  wire [511:0] _out_write_req_T_125 = _out_write_req_T_124 | _out_write_req_T_62; // @[Mux.scala 27:73]
  wire [511:0] out_write_req_data = _out_write_req_T_125 | _out_write_req_T_63; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_127 = out_write_index_0 ? mshr_0_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_128 = out_write_index_1 ? mshr_1_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_129 = out_write_index_2 ? mshr_2_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_130 = out_write_index_3 ? mshr_3_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_131 = out_write_index_4 ? mshr_4_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_132 = out_write_index_5 ? mshr_5_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_133 = out_write_index_6 ? mshr_6_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_134 = out_write_index_7 ? mshr_7_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_135 = out_write_index_8 ? mshr_8_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_136 = out_write_index_9 ? mshr_9_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_137 = out_write_index_10 ? mshr_10_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_138 = out_write_index_11 ? mshr_11_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_139 = out_write_index_12 ? mshr_12_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_140 = out_write_index_13 ? mshr_13_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_141 = out_write_index_14 ? mshr_14_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_142 = out_write_index_15 ? mshr_15_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_143 = out_write_index_16 ? mshr_16_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_144 = out_write_index_17 ? mshr_17_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_145 = out_write_index_18 ? mshr_18_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_146 = out_write_index_19 ? mshr_19_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_147 = out_write_index_20 ? mshr_20_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_148 = out_write_index_21 ? mshr_21_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_149 = out_write_index_22 ? mshr_22_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_150 = out_write_index_23 ? mshr_23_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_151 = out_write_index_24 ? mshr_24_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_152 = out_write_index_25 ? mshr_25_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_153 = out_write_index_26 ? mshr_26_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_154 = out_write_index_27 ? mshr_27_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_155 = out_write_index_28 ? mshr_28_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_156 = out_write_index_29 ? mshr_29_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_157 = out_write_index_30 ? mshr_30_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_158 = out_write_index_31 ? mshr_31_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_159 = out_write_index_32 ? mshr_32_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_160 = out_write_index_33 ? mshr_33_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_161 = out_write_index_34 ? mshr_34_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_162 = out_write_index_35 ? mshr_35_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_163 = out_write_index_36 ? mshr_36_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_164 = out_write_index_37 ? mshr_37_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_165 = out_write_index_38 ? mshr_38_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_166 = out_write_index_39 ? mshr_39_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_167 = out_write_index_40 ? mshr_40_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_168 = out_write_index_41 ? mshr_41_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_169 = out_write_index_42 ? mshr_42_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_170 = out_write_index_43 ? mshr_43_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_171 = out_write_index_44 ? mshr_44_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_172 = out_write_index_45 ? mshr_45_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_173 = out_write_index_46 ? mshr_46_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_174 = out_write_index_47 ? mshr_47_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_175 = out_write_index_48 ? mshr_48_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_176 = out_write_index_49 ? mshr_49_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_177 = out_write_index_50 ? mshr_50_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_178 = out_write_index_51 ? mshr_51_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_179 = out_write_index_52 ? mshr_52_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_180 = out_write_index_53 ? mshr_53_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_181 = out_write_index_54 ? mshr_54_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_182 = out_write_index_55 ? mshr_55_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_183 = out_write_index_56 ? mshr_56_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_184 = out_write_index_57 ? mshr_57_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_185 = out_write_index_58 ? mshr_58_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_186 = out_write_index_59 ? mshr_59_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_187 = out_write_index_60 ? mshr_60_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_188 = out_write_index_61 ? mshr_61_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_189 = out_write_index_62 ? mshr_62_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_190 = out_write_index_63 ? mshr_63_io_master_req_mask : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_191 = _out_write_req_T_127 | _out_write_req_T_128; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_192 = _out_write_req_T_191 | _out_write_req_T_129; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_193 = _out_write_req_T_192 | _out_write_req_T_130; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_194 = _out_write_req_T_193 | _out_write_req_T_131; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_195 = _out_write_req_T_194 | _out_write_req_T_132; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_196 = _out_write_req_T_195 | _out_write_req_T_133; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_197 = _out_write_req_T_196 | _out_write_req_T_134; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_198 = _out_write_req_T_197 | _out_write_req_T_135; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_199 = _out_write_req_T_198 | _out_write_req_T_136; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_200 = _out_write_req_T_199 | _out_write_req_T_137; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_201 = _out_write_req_T_200 | _out_write_req_T_138; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_202 = _out_write_req_T_201 | _out_write_req_T_139; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_203 = _out_write_req_T_202 | _out_write_req_T_140; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_204 = _out_write_req_T_203 | _out_write_req_T_141; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_205 = _out_write_req_T_204 | _out_write_req_T_142; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_206 = _out_write_req_T_205 | _out_write_req_T_143; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_207 = _out_write_req_T_206 | _out_write_req_T_144; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_208 = _out_write_req_T_207 | _out_write_req_T_145; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_209 = _out_write_req_T_208 | _out_write_req_T_146; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_210 = _out_write_req_T_209 | _out_write_req_T_147; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_211 = _out_write_req_T_210 | _out_write_req_T_148; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_212 = _out_write_req_T_211 | _out_write_req_T_149; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_213 = _out_write_req_T_212 | _out_write_req_T_150; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_214 = _out_write_req_T_213 | _out_write_req_T_151; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_215 = _out_write_req_T_214 | _out_write_req_T_152; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_216 = _out_write_req_T_215 | _out_write_req_T_153; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_217 = _out_write_req_T_216 | _out_write_req_T_154; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_218 = _out_write_req_T_217 | _out_write_req_T_155; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_219 = _out_write_req_T_218 | _out_write_req_T_156; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_220 = _out_write_req_T_219 | _out_write_req_T_157; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_221 = _out_write_req_T_220 | _out_write_req_T_158; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_222 = _out_write_req_T_221 | _out_write_req_T_159; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_223 = _out_write_req_T_222 | _out_write_req_T_160; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_224 = _out_write_req_T_223 | _out_write_req_T_161; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_225 = _out_write_req_T_224 | _out_write_req_T_162; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_226 = _out_write_req_T_225 | _out_write_req_T_163; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_227 = _out_write_req_T_226 | _out_write_req_T_164; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_228 = _out_write_req_T_227 | _out_write_req_T_165; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_229 = _out_write_req_T_228 | _out_write_req_T_166; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_230 = _out_write_req_T_229 | _out_write_req_T_167; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_231 = _out_write_req_T_230 | _out_write_req_T_168; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_232 = _out_write_req_T_231 | _out_write_req_T_169; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_233 = _out_write_req_T_232 | _out_write_req_T_170; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_234 = _out_write_req_T_233 | _out_write_req_T_171; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_235 = _out_write_req_T_234 | _out_write_req_T_172; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_236 = _out_write_req_T_235 | _out_write_req_T_173; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_237 = _out_write_req_T_236 | _out_write_req_T_174; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_238 = _out_write_req_T_237 | _out_write_req_T_175; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_239 = _out_write_req_T_238 | _out_write_req_T_176; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_240 = _out_write_req_T_239 | _out_write_req_T_177; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_241 = _out_write_req_T_240 | _out_write_req_T_178; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_242 = _out_write_req_T_241 | _out_write_req_T_179; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_243 = _out_write_req_T_242 | _out_write_req_T_180; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_244 = _out_write_req_T_243 | _out_write_req_T_181; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_245 = _out_write_req_T_244 | _out_write_req_T_182; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_246 = _out_write_req_T_245 | _out_write_req_T_183; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_247 = _out_write_req_T_246 | _out_write_req_T_184; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_248 = _out_write_req_T_247 | _out_write_req_T_185; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_249 = _out_write_req_T_248 | _out_write_req_T_186; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_250 = _out_write_req_T_249 | _out_write_req_T_187; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_251 = _out_write_req_T_250 | _out_write_req_T_188; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_252 = _out_write_req_T_251 | _out_write_req_T_189; // @[Mux.scala 27:73]
  wire [63:0] out_write_req_mask = _out_write_req_T_252 | _out_write_req_T_190; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_254 = out_write_index_0 ? mshr_0_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_255 = out_write_index_1 ? mshr_1_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_256 = out_write_index_2 ? mshr_2_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_257 = out_write_index_3 ? mshr_3_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_258 = out_write_index_4 ? mshr_4_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_259 = out_write_index_5 ? mshr_5_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_260 = out_write_index_6 ? mshr_6_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_261 = out_write_index_7 ? mshr_7_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_262 = out_write_index_8 ? mshr_8_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_263 = out_write_index_9 ? mshr_9_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_264 = out_write_index_10 ? mshr_10_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_265 = out_write_index_11 ? mshr_11_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_266 = out_write_index_12 ? mshr_12_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_267 = out_write_index_13 ? mshr_13_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_268 = out_write_index_14 ? mshr_14_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_269 = out_write_index_15 ? mshr_15_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_270 = out_write_index_16 ? mshr_16_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_271 = out_write_index_17 ? mshr_17_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_272 = out_write_index_18 ? mshr_18_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_273 = out_write_index_19 ? mshr_19_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_274 = out_write_index_20 ? mshr_20_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_275 = out_write_index_21 ? mshr_21_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_276 = out_write_index_22 ? mshr_22_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_277 = out_write_index_23 ? mshr_23_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_278 = out_write_index_24 ? mshr_24_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_279 = out_write_index_25 ? mshr_25_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_280 = out_write_index_26 ? mshr_26_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_281 = out_write_index_27 ? mshr_27_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_282 = out_write_index_28 ? mshr_28_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_283 = out_write_index_29 ? mshr_29_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_284 = out_write_index_30 ? mshr_30_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_285 = out_write_index_31 ? mshr_31_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_286 = out_write_index_32 ? mshr_32_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_287 = out_write_index_33 ? mshr_33_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_288 = out_write_index_34 ? mshr_34_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_289 = out_write_index_35 ? mshr_35_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_290 = out_write_index_36 ? mshr_36_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_291 = out_write_index_37 ? mshr_37_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_292 = out_write_index_38 ? mshr_38_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_293 = out_write_index_39 ? mshr_39_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_294 = out_write_index_40 ? mshr_40_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_295 = out_write_index_41 ? mshr_41_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_296 = out_write_index_42 ? mshr_42_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_297 = out_write_index_43 ? mshr_43_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_298 = out_write_index_44 ? mshr_44_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_299 = out_write_index_45 ? mshr_45_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_300 = out_write_index_46 ? mshr_46_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_301 = out_write_index_47 ? mshr_47_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_302 = out_write_index_48 ? mshr_48_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_303 = out_write_index_49 ? mshr_49_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_304 = out_write_index_50 ? mshr_50_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_305 = out_write_index_51 ? mshr_51_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_306 = out_write_index_52 ? mshr_52_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_307 = out_write_index_53 ? mshr_53_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_308 = out_write_index_54 ? mshr_54_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_309 = out_write_index_55 ? mshr_55_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_310 = out_write_index_56 ? mshr_56_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_311 = out_write_index_57 ? mshr_57_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_312 = out_write_index_58 ? mshr_58_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_313 = out_write_index_59 ? mshr_59_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_314 = out_write_index_60 ? mshr_60_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_315 = out_write_index_61 ? mshr_61_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_316 = out_write_index_62 ? mshr_62_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_317 = out_write_index_63 ? mshr_63_io_master_req_addr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_318 = _out_write_req_T_254 | _out_write_req_T_255; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_319 = _out_write_req_T_318 | _out_write_req_T_256; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_320 = _out_write_req_T_319 | _out_write_req_T_257; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_321 = _out_write_req_T_320 | _out_write_req_T_258; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_322 = _out_write_req_T_321 | _out_write_req_T_259; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_323 = _out_write_req_T_322 | _out_write_req_T_260; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_324 = _out_write_req_T_323 | _out_write_req_T_261; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_325 = _out_write_req_T_324 | _out_write_req_T_262; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_326 = _out_write_req_T_325 | _out_write_req_T_263; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_327 = _out_write_req_T_326 | _out_write_req_T_264; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_328 = _out_write_req_T_327 | _out_write_req_T_265; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_329 = _out_write_req_T_328 | _out_write_req_T_266; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_330 = _out_write_req_T_329 | _out_write_req_T_267; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_331 = _out_write_req_T_330 | _out_write_req_T_268; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_332 = _out_write_req_T_331 | _out_write_req_T_269; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_333 = _out_write_req_T_332 | _out_write_req_T_270; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_334 = _out_write_req_T_333 | _out_write_req_T_271; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_335 = _out_write_req_T_334 | _out_write_req_T_272; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_336 = _out_write_req_T_335 | _out_write_req_T_273; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_337 = _out_write_req_T_336 | _out_write_req_T_274; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_338 = _out_write_req_T_337 | _out_write_req_T_275; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_339 = _out_write_req_T_338 | _out_write_req_T_276; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_340 = _out_write_req_T_339 | _out_write_req_T_277; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_341 = _out_write_req_T_340 | _out_write_req_T_278; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_342 = _out_write_req_T_341 | _out_write_req_T_279; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_343 = _out_write_req_T_342 | _out_write_req_T_280; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_344 = _out_write_req_T_343 | _out_write_req_T_281; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_345 = _out_write_req_T_344 | _out_write_req_T_282; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_346 = _out_write_req_T_345 | _out_write_req_T_283; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_347 = _out_write_req_T_346 | _out_write_req_T_284; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_348 = _out_write_req_T_347 | _out_write_req_T_285; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_349 = _out_write_req_T_348 | _out_write_req_T_286; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_350 = _out_write_req_T_349 | _out_write_req_T_287; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_351 = _out_write_req_T_350 | _out_write_req_T_288; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_352 = _out_write_req_T_351 | _out_write_req_T_289; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_353 = _out_write_req_T_352 | _out_write_req_T_290; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_354 = _out_write_req_T_353 | _out_write_req_T_291; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_355 = _out_write_req_T_354 | _out_write_req_T_292; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_356 = _out_write_req_T_355 | _out_write_req_T_293; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_357 = _out_write_req_T_356 | _out_write_req_T_294; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_358 = _out_write_req_T_357 | _out_write_req_T_295; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_359 = _out_write_req_T_358 | _out_write_req_T_296; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_360 = _out_write_req_T_359 | _out_write_req_T_297; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_361 = _out_write_req_T_360 | _out_write_req_T_298; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_362 = _out_write_req_T_361 | _out_write_req_T_299; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_363 = _out_write_req_T_362 | _out_write_req_T_300; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_364 = _out_write_req_T_363 | _out_write_req_T_301; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_365 = _out_write_req_T_364 | _out_write_req_T_302; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_366 = _out_write_req_T_365 | _out_write_req_T_303; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_367 = _out_write_req_T_366 | _out_write_req_T_304; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_368 = _out_write_req_T_367 | _out_write_req_T_305; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_369 = _out_write_req_T_368 | _out_write_req_T_306; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_370 = _out_write_req_T_369 | _out_write_req_T_307; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_371 = _out_write_req_T_370 | _out_write_req_T_308; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_372 = _out_write_req_T_371 | _out_write_req_T_309; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_373 = _out_write_req_T_372 | _out_write_req_T_310; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_374 = _out_write_req_T_373 | _out_write_req_T_311; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_375 = _out_write_req_T_374 | _out_write_req_T_312; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_376 = _out_write_req_T_375 | _out_write_req_T_313; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_377 = _out_write_req_T_376 | _out_write_req_T_314; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_378 = _out_write_req_T_377 | _out_write_req_T_315; // @[Mux.scala 27:73]
  wire [63:0] _out_write_req_T_379 = _out_write_req_T_378 | _out_write_req_T_316; // @[Mux.scala 27:73]
  wire [63:0] out_write_req_addr = _out_write_req_T_379 | _out_write_req_T_317; // @[Mux.scala 27:73]
  wire [7:0] bundleOut_0_awvalid_lo_lo_lo = {has_write_req_7,has_write_req_6,has_write_req_5,has_write_req_4,
    has_write_req_3,has_write_req_2,has_write_req_1,has_write_req_0}; // @[AXI4FakeDMA.scala 199:35]
  wire [15:0] bundleOut_0_awvalid_lo_lo = {has_write_req_15,has_write_req_14,has_write_req_13,has_write_req_12,
    has_write_req_11,has_write_req_10,has_write_req_9,has_write_req_8,bundleOut_0_awvalid_lo_lo_lo}; // @[AXI4FakeDMA.scala 199:35]
  wire [7:0] bundleOut_0_awvalid_lo_hi_lo = {has_write_req_23,has_write_req_22,has_write_req_21,has_write_req_20,
    has_write_req_19,has_write_req_18,has_write_req_17,has_write_req_16}; // @[AXI4FakeDMA.scala 199:35]
  wire [31:0] bundleOut_0_awvalid_lo = {has_write_req_31,has_write_req_30,has_write_req_29,has_write_req_28,
    has_write_req_27,has_write_req_26,has_write_req_25,has_write_req_24,bundleOut_0_awvalid_lo_hi_lo,
    bundleOut_0_awvalid_lo_lo}; // @[AXI4FakeDMA.scala 199:35]
  wire [7:0] bundleOut_0_awvalid_hi_lo_lo = {has_write_req_39,has_write_req_38,has_write_req_37,has_write_req_36,
    has_write_req_35,has_write_req_34,has_write_req_33,has_write_req_32}; // @[AXI4FakeDMA.scala 199:35]
  wire [15:0] bundleOut_0_awvalid_hi_lo = {has_write_req_47,has_write_req_46,has_write_req_45,has_write_req_44,
    has_write_req_43,has_write_req_42,has_write_req_41,has_write_req_40,bundleOut_0_awvalid_hi_lo_lo}; // @[AXI4FakeDMA.scala 199:35]
  wire [7:0] bundleOut_0_awvalid_hi_hi_lo = {has_write_req_55,has_write_req_54,has_write_req_53,has_write_req_52,
    has_write_req_51,has_write_req_50,has_write_req_49,has_write_req_48}; // @[AXI4FakeDMA.scala 199:35]
  wire [31:0] bundleOut_0_awvalid_hi = {has_write_req_63,has_write_req_62,has_write_req_61,has_write_req_60,
    has_write_req_59,has_write_req_58,has_write_req_57,has_write_req_56,bundleOut_0_awvalid_hi_hi_lo,
    bundleOut_0_awvalid_hi_lo}; // @[AXI4FakeDMA.scala 199:35]
  wire [63:0] _bundleOut_0_awvalid_T = {bundleOut_0_awvalid_hi,bundleOut_0_awvalid_lo}; // @[AXI4FakeDMA.scala 199:35]
  wire [7:0] bundleOut_0_awid_lo_lo_lo = {out_write_index_7,out_write_index_6,out_write_index_5,out_write_index_4,
    out_write_index_3,out_write_index_2,out_write_index_1,out_write_index_0}; // @[Cat.scala 31:58]
  wire [15:0] bundleOut_0_awid_lo_lo = {out_write_index_15,out_write_index_14,out_write_index_13,
    out_write_index_12,out_write_index_11,out_write_index_10,out_write_index_9,out_write_index_8,
    bundleOut_0_awid_lo_lo_lo}; // @[Cat.scala 31:58]
  wire [7:0] bundleOut_0_awid_lo_hi_lo = {out_write_index_23,out_write_index_22,out_write_index_21,
    out_write_index_20,out_write_index_19,out_write_index_18,out_write_index_17,out_write_index_16}; // @[Cat.scala 31:58]
  wire [31:0] bundleOut_0_awid_lo = {out_write_index_31,out_write_index_30,out_write_index_29,out_write_index_28,
    out_write_index_27,out_write_index_26,out_write_index_25,out_write_index_24,bundleOut_0_awid_lo_hi_lo,
    bundleOut_0_awid_lo_lo}; // @[Cat.scala 31:58]
  wire [7:0] bundleOut_0_awid_hi_lo_lo = {out_write_index_39,out_write_index_38,out_write_index_37,
    out_write_index_36,out_write_index_35,out_write_index_34,out_write_index_33,out_write_index_32}; // @[Cat.scala 31:58]
  wire [15:0] bundleOut_0_awid_hi_lo = {out_write_index_47,out_write_index_46,out_write_index_45,
    out_write_index_44,out_write_index_43,out_write_index_42,out_write_index_41,out_write_index_40,
    bundleOut_0_awid_hi_lo_lo}; // @[Cat.scala 31:58]
  wire [7:0] bundleOut_0_awid_hi_hi_lo = {out_write_index_55,out_write_index_54,out_write_index_53,
    out_write_index_52,out_write_index_51,out_write_index_50,out_write_index_49,out_write_index_48}; // @[Cat.scala 31:58]
  wire [31:0] bundleOut_0_awid_hi = {out_write_index_63,out_write_index_62,out_write_index_61,out_write_index_60,
    out_write_index_59,out_write_index_58,out_write_index_57,out_write_index_56,bundleOut_0_awid_hi_hi_lo,
    bundleOut_0_awid_hi_lo}; // @[Cat.scala 31:58]
  wire [63:0] _bundleOut_0_awid_T = {bundleOut_0_awid_hi,bundleOut_0_awid_lo}; // @[Cat.scala 31:58]
  wire [31:0] bundleOut_0_awid_hi_1 = _bundleOut_0_awid_T[63:32]; // @[OneHot.scala 30:18]
  wire [31:0] bundleOut_0_awid_lo_1 = _bundleOut_0_awid_T[31:0]; // @[OneHot.scala 31:18]
  wire  _bundleOut_0_awid_T_1 = |bundleOut_0_awid_hi_1; // @[OneHot.scala 32:14]
  wire [31:0] _bundleOut_0_awid_T_2 = bundleOut_0_awid_hi_1 | bundleOut_0_awid_lo_1; // @[OneHot.scala 32:28]
  wire [15:0] bundleOut_0_awid_hi_2 = _bundleOut_0_awid_T_2[31:16]; // @[OneHot.scala 30:18]
  wire [15:0] bundleOut_0_awid_lo_2 = _bundleOut_0_awid_T_2[15:0]; // @[OneHot.scala 31:18]
  wire  _bundleOut_0_awid_T_3 = |bundleOut_0_awid_hi_2; // @[OneHot.scala 32:14]
  wire [15:0] _bundleOut_0_awid_T_4 = bundleOut_0_awid_hi_2 | bundleOut_0_awid_lo_2; // @[OneHot.scala 32:28]
  wire [7:0] bundleOut_0_awid_hi_3 = _bundleOut_0_awid_T_4[15:8]; // @[OneHot.scala 30:18]
  wire [7:0] bundleOut_0_awid_lo_3 = _bundleOut_0_awid_T_4[7:0]; // @[OneHot.scala 31:18]
  wire  _bundleOut_0_awid_T_5 = |bundleOut_0_awid_hi_3; // @[OneHot.scala 32:14]
  wire [7:0] _bundleOut_0_awid_T_6 = bundleOut_0_awid_hi_3 | bundleOut_0_awid_lo_3; // @[OneHot.scala 32:28]
  wire [3:0] bundleOut_0_awid_hi_4 = _bundleOut_0_awid_T_6[7:4]; // @[OneHot.scala 30:18]
  wire [3:0] bundleOut_0_awid_lo_4 = _bundleOut_0_awid_T_6[3:0]; // @[OneHot.scala 31:18]
  wire  _bundleOut_0_awid_T_7 = |bundleOut_0_awid_hi_4; // @[OneHot.scala 32:14]
  wire [3:0] _bundleOut_0_awid_T_8 = bundleOut_0_awid_hi_4 | bundleOut_0_awid_lo_4; // @[OneHot.scala 32:28]
  wire [1:0] bundleOut_0_awid_hi_5 = _bundleOut_0_awid_T_8[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] bundleOut_0_awid_lo_5 = _bundleOut_0_awid_T_8[1:0]; // @[OneHot.scala 31:18]
  wire  _bundleOut_0_awid_T_9 = |bundleOut_0_awid_hi_5; // @[OneHot.scala 32:14]
  wire [1:0] _bundleOut_0_awid_T_10 = bundleOut_0_awid_hi_5 | bundleOut_0_awid_lo_5; // @[OneHot.scala 32:28]
  wire [5:0] _bundleOut_0_awid_T_16 = {_bundleOut_0_awid_T_1,_bundleOut_0_awid_T_3,
    _bundleOut_0_awid_T_5,_bundleOut_0_awid_T_7,_bundleOut_0_awid_T_9,_bundleOut_0_awid_T_10[1]}
    ; // @[Cat.scala 31:58]
  wire  _read_fire_T = auto_dma_out_arready & out_arvalid; // @[Decoupled.scala 50:35]
  wire  read_fire = _read_fire_T & out_read_index_0; // @[AXI4FakeDMA.scala 209:35]
  reg  w_valid; // @[AXI4FakeDMA.scala 215:26]
  wire  out_awvalid = w_valid ? 1'h0 : |_bundleOut_0_awvalid_T; // @[AXI4FakeDMA.scala 199:18 222:20 223:20]
  wire  _write_fire_T = auto_dma_out_awready & out_awvalid; // @[Decoupled.scala 50:35]
  wire  write_fire = _write_fire_T & out_write_index_0; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_1 = _read_fire_T & out_read_index_1; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_1 = _write_fire_T & out_write_index_1; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_2 = _read_fire_T & out_read_index_2; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_2 = _write_fire_T & out_write_index_2; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_3 = _read_fire_T & out_read_index_3; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_3 = _write_fire_T & out_write_index_3; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_4 = _read_fire_T & out_read_index_4; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_4 = _write_fire_T & out_write_index_4; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_5 = _read_fire_T & out_read_index_5; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_5 = _write_fire_T & out_write_index_5; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_6 = _read_fire_T & out_read_index_6; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_6 = _write_fire_T & out_write_index_6; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_7 = _read_fire_T & out_read_index_7; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_7 = _write_fire_T & out_write_index_7; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_8 = _read_fire_T & out_read_index_8; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_8 = _write_fire_T & out_write_index_8; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_9 = _read_fire_T & out_read_index_9; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_9 = _write_fire_T & out_write_index_9; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_10 = _read_fire_T & out_read_index_10; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_10 = _write_fire_T & out_write_index_10; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_11 = _read_fire_T & out_read_index_11; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_11 = _write_fire_T & out_write_index_11; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_12 = _read_fire_T & out_read_index_12; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_12 = _write_fire_T & out_write_index_12; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_13 = _read_fire_T & out_read_index_13; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_13 = _write_fire_T & out_write_index_13; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_14 = _read_fire_T & out_read_index_14; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_14 = _write_fire_T & out_write_index_14; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_15 = _read_fire_T & out_read_index_15; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_15 = _write_fire_T & out_write_index_15; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_16 = _read_fire_T & out_read_index_16; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_16 = _write_fire_T & out_write_index_16; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_17 = _read_fire_T & out_read_index_17; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_17 = _write_fire_T & out_write_index_17; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_18 = _read_fire_T & out_read_index_18; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_18 = _write_fire_T & out_write_index_18; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_19 = _read_fire_T & out_read_index_19; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_19 = _write_fire_T & out_write_index_19; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_20 = _read_fire_T & out_read_index_20; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_20 = _write_fire_T & out_write_index_20; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_21 = _read_fire_T & out_read_index_21; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_21 = _write_fire_T & out_write_index_21; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_22 = _read_fire_T & out_read_index_22; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_22 = _write_fire_T & out_write_index_22; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_23 = _read_fire_T & out_read_index_23; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_23 = _write_fire_T & out_write_index_23; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_24 = _read_fire_T & out_read_index_24; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_24 = _write_fire_T & out_write_index_24; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_25 = _read_fire_T & out_read_index_25; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_25 = _write_fire_T & out_write_index_25; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_26 = _read_fire_T & out_read_index_26; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_26 = _write_fire_T & out_write_index_26; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_27 = _read_fire_T & out_read_index_27; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_27 = _write_fire_T & out_write_index_27; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_28 = _read_fire_T & out_read_index_28; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_28 = _write_fire_T & out_write_index_28; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_29 = _read_fire_T & out_read_index_29; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_29 = _write_fire_T & out_write_index_29; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_30 = _read_fire_T & out_read_index_30; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_30 = _write_fire_T & out_write_index_30; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_31 = _read_fire_T & out_read_index_31; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_31 = _write_fire_T & out_write_index_31; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_32 = _read_fire_T & out_read_index_32; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_32 = _write_fire_T & out_write_index_32; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_33 = _read_fire_T & out_read_index_33; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_33 = _write_fire_T & out_write_index_33; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_34 = _read_fire_T & out_read_index_34; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_34 = _write_fire_T & out_write_index_34; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_35 = _read_fire_T & out_read_index_35; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_35 = _write_fire_T & out_write_index_35; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_36 = _read_fire_T & out_read_index_36; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_36 = _write_fire_T & out_write_index_36; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_37 = _read_fire_T & out_read_index_37; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_37 = _write_fire_T & out_write_index_37; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_38 = _read_fire_T & out_read_index_38; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_38 = _write_fire_T & out_write_index_38; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_39 = _read_fire_T & out_read_index_39; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_39 = _write_fire_T & out_write_index_39; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_40 = _read_fire_T & out_read_index_40; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_40 = _write_fire_T & out_write_index_40; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_41 = _read_fire_T & out_read_index_41; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_41 = _write_fire_T & out_write_index_41; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_42 = _read_fire_T & out_read_index_42; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_42 = _write_fire_T & out_write_index_42; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_43 = _read_fire_T & out_read_index_43; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_43 = _write_fire_T & out_write_index_43; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_44 = _read_fire_T & out_read_index_44; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_44 = _write_fire_T & out_write_index_44; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_45 = _read_fire_T & out_read_index_45; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_45 = _write_fire_T & out_write_index_45; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_46 = _read_fire_T & out_read_index_46; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_46 = _write_fire_T & out_write_index_46; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_47 = _read_fire_T & out_read_index_47; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_47 = _write_fire_T & out_write_index_47; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_48 = _read_fire_T & out_read_index_48; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_48 = _write_fire_T & out_write_index_48; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_49 = _read_fire_T & out_read_index_49; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_49 = _write_fire_T & out_write_index_49; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_50 = _read_fire_T & out_read_index_50; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_50 = _write_fire_T & out_write_index_50; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_51 = _read_fire_T & out_read_index_51; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_51 = _write_fire_T & out_write_index_51; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_52 = _read_fire_T & out_read_index_52; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_52 = _write_fire_T & out_write_index_52; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_53 = _read_fire_T & out_read_index_53; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_53 = _write_fire_T & out_write_index_53; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_54 = _read_fire_T & out_read_index_54; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_54 = _write_fire_T & out_write_index_54; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_55 = _read_fire_T & out_read_index_55; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_55 = _write_fire_T & out_write_index_55; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_56 = _read_fire_T & out_read_index_56; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_56 = _write_fire_T & out_write_index_56; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_57 = _read_fire_T & out_read_index_57; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_57 = _write_fire_T & out_write_index_57; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_58 = _read_fire_T & out_read_index_58; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_58 = _write_fire_T & out_write_index_58; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_59 = _read_fire_T & out_read_index_59; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_59 = _write_fire_T & out_write_index_59; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_60 = _read_fire_T & out_read_index_60; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_60 = _write_fire_T & out_write_index_60; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_61 = _read_fire_T & out_read_index_61; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_61 = _write_fire_T & out_write_index_61; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_62 = _read_fire_T & out_read_index_62; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_62 = _write_fire_T & out_write_index_62; // @[AXI4FakeDMA.scala 210:36]
  wire  read_fire_63 = _read_fire_T & out_read_index_63; // @[AXI4FakeDMA.scala 209:35]
  wire  write_fire_63 = _write_fire_T & out_write_index_63; // @[AXI4FakeDMA.scala 210:36]
  wire  _T_495 = auto_dma_out_wready & w_valid; // @[Decoupled.scala 50:35]
  reg  beatCount; // @[AXI4FakeDMA.scala 225:28]
  wire  _GEN_275 = _T_495 & beatCount ? 1'h0 : w_valid; // @[AXI4FakeDMA.scala 218:47 219:15 215:26]
  wire  _GEN_276 = _write_fire_T | _GEN_275; // @[AXI4FakeDMA.scala 216:24 217:15]
  reg [63:0] w_mask; // @[Reg.scala 16:16]
  reg [511:0] w_data; // @[Reg.scala 16:16]
  wire  read_resp_fire = auto_dma_out_rvalid & auto_dma_out_rid == 8'h0; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire = auto_dma_out_bvalid & auto_dma_out_bid == 8'h0; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_1 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h1; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_1 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h1; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_2 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h2; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_2 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h2; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_3 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h3; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_3 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h3; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_4 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h4; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_4 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h4; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_5 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h5; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_5 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h5; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_6 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h6; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_6 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h6; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_7 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h7; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_7 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h7; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_8 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h8; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_8 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h8; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_9 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h9; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_9 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h9; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_10 = auto_dma_out_rvalid & auto_dma_out_rid == 8'ha; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_10 = auto_dma_out_bvalid & auto_dma_out_bid == 8'ha; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_11 = auto_dma_out_rvalid & auto_dma_out_rid == 8'hb; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_11 = auto_dma_out_bvalid & auto_dma_out_bid == 8'hb; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_12 = auto_dma_out_rvalid & auto_dma_out_rid == 8'hc; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_12 = auto_dma_out_bvalid & auto_dma_out_bid == 8'hc; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_13 = auto_dma_out_rvalid & auto_dma_out_rid == 8'hd; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_13 = auto_dma_out_bvalid & auto_dma_out_bid == 8'hd; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_14 = auto_dma_out_rvalid & auto_dma_out_rid == 8'he; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_14 = auto_dma_out_bvalid & auto_dma_out_bid == 8'he; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_15 = auto_dma_out_rvalid & auto_dma_out_rid == 8'hf; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_15 = auto_dma_out_bvalid & auto_dma_out_bid == 8'hf; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_16 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h10; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_16 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h10; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_17 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h11; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_17 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h11; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_18 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h12; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_18 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h12; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_19 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h13; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_19 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h13; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_20 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h14; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_20 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h14; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_21 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h15; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_21 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h15; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_22 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h16; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_22 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h16; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_23 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h17; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_23 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h17; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_24 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h18; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_24 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h18; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_25 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h19; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_25 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h19; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_26 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h1a; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_26 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h1a; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_27 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h1b; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_27 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h1b; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_28 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h1c; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_28 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h1c; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_29 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h1d; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_29 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h1d; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_30 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h1e; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_30 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h1e; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_31 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h1f; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_31 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h1f; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_32 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h20; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_32 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h20; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_33 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h21; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_33 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h21; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_34 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h22; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_34 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h22; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_35 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h23; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_35 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h23; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_36 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h24; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_36 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h24; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_37 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h25; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_37 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h25; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_38 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h26; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_38 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h26; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_39 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h27; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_39 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h27; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_40 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h28; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_40 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h28; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_41 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h29; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_41 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h29; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_42 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h2a; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_42 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h2a; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_43 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h2b; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_43 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h2b; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_44 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h2c; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_44 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h2c; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_45 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h2d; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_45 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h2d; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_46 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h2e; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_46 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h2e; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_47 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h2f; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_47 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h2f; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_48 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h30; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_48 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h30; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_49 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h31; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_49 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h31; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_50 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h32; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_50 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h32; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_51 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h33; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_51 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h33; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_52 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h34; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_52 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h34; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_53 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h35; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_53 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h35; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_54 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h36; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_54 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h36; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_55 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h37; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_55 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h37; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_56 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h38; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_56 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h38; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_57 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h39; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_57 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h39; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_58 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h3a; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_58 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h3a; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_59 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h3b; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_59 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h3b; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_60 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h3c; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_60 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h3c; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_61 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h3d; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_61 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h3d; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_62 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h3e; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_62 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h3e; // @[AXI4FakeDMA.scala 242:40]
  wire  read_resp_fire_63 = auto_dma_out_rvalid & auto_dma_out_rid == 8'h3f; // @[AXI4FakeDMA.scala 241:39]
  wire  write_resp_fire_63 = auto_dma_out_bvalid & auto_dma_out_bid == 8'h3f; // @[AXI4FakeDMA.scala 242:40]
  wire [7:0] in_awlen = auto_in_awlen; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  wire [2:0] in_awsize = auto_in_awsize; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  wire  in_awlock = auto_in_awlock; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  wire [3:0] in_awcache = auto_in_awcache; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  wire [2:0] in_awprot = auto_in_awprot; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  wire [3:0] in_awqos = auto_in_awqos; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  wire  in_bid = bundleIn_0_bid_r; // @[Nodes.scala 1210:84 AXI4SlaveModule.scala 177:16]
  wire [1:0] in_bresp = 2'h0; // @[Nodes.scala 1210:84 AXI4SlaveModule.scala 174:18]
  wire [2:0] in_arsize = auto_in_arsize; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  wire  in_arlock = auto_in_arlock; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  wire [3:0] in_arcache = auto_in_arcache; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  wire [2:0] in_arprot = auto_in_arprot; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  wire [3:0] in_arqos = auto_in_arqos; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  wire  in_rid = bundleIn_0_rid_r; // @[Nodes.scala 1210:84 AXI4SlaveModule.scala 179:16]
  wire [63:0] in_rdata = _GEN_10[13] ? enable : _GEN_81; // @[AXI4FakeDMA.scala 158:26]
  wire [1:0] in_rresp = 2'h0; // @[Nodes.scala 1210:84 AXI4SlaveModule.scala 154:18]
  DMAFakeMSHR mshr_0 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_0_clock),
    .reset(mshr_0_reset),
    .io_enable(mshr_0_io_enable),
    .io_slave_wen(mshr_0_io_slave_wen),
    .io_slave_addr(mshr_0_io_slave_addr),
    .io_slave_rdata(mshr_0_io_slave_rdata),
    .io_slave_wdata(mshr_0_io_slave_wdata),
    .io_master_req_valid(mshr_0_io_master_req_valid),
    .io_master_req_ready(mshr_0_io_master_req_ready),
    .io_master_req_is_write(mshr_0_io_master_req_is_write),
    .io_master_req_addr(mshr_0_io_master_req_addr),
    .io_master_req_mask(mshr_0_io_master_req_mask),
    .io_master_req_data(mshr_0_io_master_req_data),
    .io_master_resp_valid(mshr_0_io_master_resp_valid),
    .io_master_resp_bits(mshr_0_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_1 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_1_clock),
    .reset(mshr_1_reset),
    .io_enable(mshr_1_io_enable),
    .io_slave_wen(mshr_1_io_slave_wen),
    .io_slave_addr(mshr_1_io_slave_addr),
    .io_slave_rdata(mshr_1_io_slave_rdata),
    .io_slave_wdata(mshr_1_io_slave_wdata),
    .io_master_req_valid(mshr_1_io_master_req_valid),
    .io_master_req_ready(mshr_1_io_master_req_ready),
    .io_master_req_is_write(mshr_1_io_master_req_is_write),
    .io_master_req_addr(mshr_1_io_master_req_addr),
    .io_master_req_mask(mshr_1_io_master_req_mask),
    .io_master_req_data(mshr_1_io_master_req_data),
    .io_master_resp_valid(mshr_1_io_master_resp_valid),
    .io_master_resp_bits(mshr_1_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_2 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_2_clock),
    .reset(mshr_2_reset),
    .io_enable(mshr_2_io_enable),
    .io_slave_wen(mshr_2_io_slave_wen),
    .io_slave_addr(mshr_2_io_slave_addr),
    .io_slave_rdata(mshr_2_io_slave_rdata),
    .io_slave_wdata(mshr_2_io_slave_wdata),
    .io_master_req_valid(mshr_2_io_master_req_valid),
    .io_master_req_ready(mshr_2_io_master_req_ready),
    .io_master_req_is_write(mshr_2_io_master_req_is_write),
    .io_master_req_addr(mshr_2_io_master_req_addr),
    .io_master_req_mask(mshr_2_io_master_req_mask),
    .io_master_req_data(mshr_2_io_master_req_data),
    .io_master_resp_valid(mshr_2_io_master_resp_valid),
    .io_master_resp_bits(mshr_2_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_3 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_3_clock),
    .reset(mshr_3_reset),
    .io_enable(mshr_3_io_enable),
    .io_slave_wen(mshr_3_io_slave_wen),
    .io_slave_addr(mshr_3_io_slave_addr),
    .io_slave_rdata(mshr_3_io_slave_rdata),
    .io_slave_wdata(mshr_3_io_slave_wdata),
    .io_master_req_valid(mshr_3_io_master_req_valid),
    .io_master_req_ready(mshr_3_io_master_req_ready),
    .io_master_req_is_write(mshr_3_io_master_req_is_write),
    .io_master_req_addr(mshr_3_io_master_req_addr),
    .io_master_req_mask(mshr_3_io_master_req_mask),
    .io_master_req_data(mshr_3_io_master_req_data),
    .io_master_resp_valid(mshr_3_io_master_resp_valid),
    .io_master_resp_bits(mshr_3_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_4 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_4_clock),
    .reset(mshr_4_reset),
    .io_enable(mshr_4_io_enable),
    .io_slave_wen(mshr_4_io_slave_wen),
    .io_slave_addr(mshr_4_io_slave_addr),
    .io_slave_rdata(mshr_4_io_slave_rdata),
    .io_slave_wdata(mshr_4_io_slave_wdata),
    .io_master_req_valid(mshr_4_io_master_req_valid),
    .io_master_req_ready(mshr_4_io_master_req_ready),
    .io_master_req_is_write(mshr_4_io_master_req_is_write),
    .io_master_req_addr(mshr_4_io_master_req_addr),
    .io_master_req_mask(mshr_4_io_master_req_mask),
    .io_master_req_data(mshr_4_io_master_req_data),
    .io_master_resp_valid(mshr_4_io_master_resp_valid),
    .io_master_resp_bits(mshr_4_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_5 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_5_clock),
    .reset(mshr_5_reset),
    .io_enable(mshr_5_io_enable),
    .io_slave_wen(mshr_5_io_slave_wen),
    .io_slave_addr(mshr_5_io_slave_addr),
    .io_slave_rdata(mshr_5_io_slave_rdata),
    .io_slave_wdata(mshr_5_io_slave_wdata),
    .io_master_req_valid(mshr_5_io_master_req_valid),
    .io_master_req_ready(mshr_5_io_master_req_ready),
    .io_master_req_is_write(mshr_5_io_master_req_is_write),
    .io_master_req_addr(mshr_5_io_master_req_addr),
    .io_master_req_mask(mshr_5_io_master_req_mask),
    .io_master_req_data(mshr_5_io_master_req_data),
    .io_master_resp_valid(mshr_5_io_master_resp_valid),
    .io_master_resp_bits(mshr_5_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_6 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_6_clock),
    .reset(mshr_6_reset),
    .io_enable(mshr_6_io_enable),
    .io_slave_wen(mshr_6_io_slave_wen),
    .io_slave_addr(mshr_6_io_slave_addr),
    .io_slave_rdata(mshr_6_io_slave_rdata),
    .io_slave_wdata(mshr_6_io_slave_wdata),
    .io_master_req_valid(mshr_6_io_master_req_valid),
    .io_master_req_ready(mshr_6_io_master_req_ready),
    .io_master_req_is_write(mshr_6_io_master_req_is_write),
    .io_master_req_addr(mshr_6_io_master_req_addr),
    .io_master_req_mask(mshr_6_io_master_req_mask),
    .io_master_req_data(mshr_6_io_master_req_data),
    .io_master_resp_valid(mshr_6_io_master_resp_valid),
    .io_master_resp_bits(mshr_6_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_7 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_7_clock),
    .reset(mshr_7_reset),
    .io_enable(mshr_7_io_enable),
    .io_slave_wen(mshr_7_io_slave_wen),
    .io_slave_addr(mshr_7_io_slave_addr),
    .io_slave_rdata(mshr_7_io_slave_rdata),
    .io_slave_wdata(mshr_7_io_slave_wdata),
    .io_master_req_valid(mshr_7_io_master_req_valid),
    .io_master_req_ready(mshr_7_io_master_req_ready),
    .io_master_req_is_write(mshr_7_io_master_req_is_write),
    .io_master_req_addr(mshr_7_io_master_req_addr),
    .io_master_req_mask(mshr_7_io_master_req_mask),
    .io_master_req_data(mshr_7_io_master_req_data),
    .io_master_resp_valid(mshr_7_io_master_resp_valid),
    .io_master_resp_bits(mshr_7_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_8 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_8_clock),
    .reset(mshr_8_reset),
    .io_enable(mshr_8_io_enable),
    .io_slave_wen(mshr_8_io_slave_wen),
    .io_slave_addr(mshr_8_io_slave_addr),
    .io_slave_rdata(mshr_8_io_slave_rdata),
    .io_slave_wdata(mshr_8_io_slave_wdata),
    .io_master_req_valid(mshr_8_io_master_req_valid),
    .io_master_req_ready(mshr_8_io_master_req_ready),
    .io_master_req_is_write(mshr_8_io_master_req_is_write),
    .io_master_req_addr(mshr_8_io_master_req_addr),
    .io_master_req_mask(mshr_8_io_master_req_mask),
    .io_master_req_data(mshr_8_io_master_req_data),
    .io_master_resp_valid(mshr_8_io_master_resp_valid),
    .io_master_resp_bits(mshr_8_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_9 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_9_clock),
    .reset(mshr_9_reset),
    .io_enable(mshr_9_io_enable),
    .io_slave_wen(mshr_9_io_slave_wen),
    .io_slave_addr(mshr_9_io_slave_addr),
    .io_slave_rdata(mshr_9_io_slave_rdata),
    .io_slave_wdata(mshr_9_io_slave_wdata),
    .io_master_req_valid(mshr_9_io_master_req_valid),
    .io_master_req_ready(mshr_9_io_master_req_ready),
    .io_master_req_is_write(mshr_9_io_master_req_is_write),
    .io_master_req_addr(mshr_9_io_master_req_addr),
    .io_master_req_mask(mshr_9_io_master_req_mask),
    .io_master_req_data(mshr_9_io_master_req_data),
    .io_master_resp_valid(mshr_9_io_master_resp_valid),
    .io_master_resp_bits(mshr_9_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_10 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_10_clock),
    .reset(mshr_10_reset),
    .io_enable(mshr_10_io_enable),
    .io_slave_wen(mshr_10_io_slave_wen),
    .io_slave_addr(mshr_10_io_slave_addr),
    .io_slave_rdata(mshr_10_io_slave_rdata),
    .io_slave_wdata(mshr_10_io_slave_wdata),
    .io_master_req_valid(mshr_10_io_master_req_valid),
    .io_master_req_ready(mshr_10_io_master_req_ready),
    .io_master_req_is_write(mshr_10_io_master_req_is_write),
    .io_master_req_addr(mshr_10_io_master_req_addr),
    .io_master_req_mask(mshr_10_io_master_req_mask),
    .io_master_req_data(mshr_10_io_master_req_data),
    .io_master_resp_valid(mshr_10_io_master_resp_valid),
    .io_master_resp_bits(mshr_10_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_11 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_11_clock),
    .reset(mshr_11_reset),
    .io_enable(mshr_11_io_enable),
    .io_slave_wen(mshr_11_io_slave_wen),
    .io_slave_addr(mshr_11_io_slave_addr),
    .io_slave_rdata(mshr_11_io_slave_rdata),
    .io_slave_wdata(mshr_11_io_slave_wdata),
    .io_master_req_valid(mshr_11_io_master_req_valid),
    .io_master_req_ready(mshr_11_io_master_req_ready),
    .io_master_req_is_write(mshr_11_io_master_req_is_write),
    .io_master_req_addr(mshr_11_io_master_req_addr),
    .io_master_req_mask(mshr_11_io_master_req_mask),
    .io_master_req_data(mshr_11_io_master_req_data),
    .io_master_resp_valid(mshr_11_io_master_resp_valid),
    .io_master_resp_bits(mshr_11_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_12 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_12_clock),
    .reset(mshr_12_reset),
    .io_enable(mshr_12_io_enable),
    .io_slave_wen(mshr_12_io_slave_wen),
    .io_slave_addr(mshr_12_io_slave_addr),
    .io_slave_rdata(mshr_12_io_slave_rdata),
    .io_slave_wdata(mshr_12_io_slave_wdata),
    .io_master_req_valid(mshr_12_io_master_req_valid),
    .io_master_req_ready(mshr_12_io_master_req_ready),
    .io_master_req_is_write(mshr_12_io_master_req_is_write),
    .io_master_req_addr(mshr_12_io_master_req_addr),
    .io_master_req_mask(mshr_12_io_master_req_mask),
    .io_master_req_data(mshr_12_io_master_req_data),
    .io_master_resp_valid(mshr_12_io_master_resp_valid),
    .io_master_resp_bits(mshr_12_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_13 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_13_clock),
    .reset(mshr_13_reset),
    .io_enable(mshr_13_io_enable),
    .io_slave_wen(mshr_13_io_slave_wen),
    .io_slave_addr(mshr_13_io_slave_addr),
    .io_slave_rdata(mshr_13_io_slave_rdata),
    .io_slave_wdata(mshr_13_io_slave_wdata),
    .io_master_req_valid(mshr_13_io_master_req_valid),
    .io_master_req_ready(mshr_13_io_master_req_ready),
    .io_master_req_is_write(mshr_13_io_master_req_is_write),
    .io_master_req_addr(mshr_13_io_master_req_addr),
    .io_master_req_mask(mshr_13_io_master_req_mask),
    .io_master_req_data(mshr_13_io_master_req_data),
    .io_master_resp_valid(mshr_13_io_master_resp_valid),
    .io_master_resp_bits(mshr_13_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_14 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_14_clock),
    .reset(mshr_14_reset),
    .io_enable(mshr_14_io_enable),
    .io_slave_wen(mshr_14_io_slave_wen),
    .io_slave_addr(mshr_14_io_slave_addr),
    .io_slave_rdata(mshr_14_io_slave_rdata),
    .io_slave_wdata(mshr_14_io_slave_wdata),
    .io_master_req_valid(mshr_14_io_master_req_valid),
    .io_master_req_ready(mshr_14_io_master_req_ready),
    .io_master_req_is_write(mshr_14_io_master_req_is_write),
    .io_master_req_addr(mshr_14_io_master_req_addr),
    .io_master_req_mask(mshr_14_io_master_req_mask),
    .io_master_req_data(mshr_14_io_master_req_data),
    .io_master_resp_valid(mshr_14_io_master_resp_valid),
    .io_master_resp_bits(mshr_14_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_15 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_15_clock),
    .reset(mshr_15_reset),
    .io_enable(mshr_15_io_enable),
    .io_slave_wen(mshr_15_io_slave_wen),
    .io_slave_addr(mshr_15_io_slave_addr),
    .io_slave_rdata(mshr_15_io_slave_rdata),
    .io_slave_wdata(mshr_15_io_slave_wdata),
    .io_master_req_valid(mshr_15_io_master_req_valid),
    .io_master_req_ready(mshr_15_io_master_req_ready),
    .io_master_req_is_write(mshr_15_io_master_req_is_write),
    .io_master_req_addr(mshr_15_io_master_req_addr),
    .io_master_req_mask(mshr_15_io_master_req_mask),
    .io_master_req_data(mshr_15_io_master_req_data),
    .io_master_resp_valid(mshr_15_io_master_resp_valid),
    .io_master_resp_bits(mshr_15_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_16 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_16_clock),
    .reset(mshr_16_reset),
    .io_enable(mshr_16_io_enable),
    .io_slave_wen(mshr_16_io_slave_wen),
    .io_slave_addr(mshr_16_io_slave_addr),
    .io_slave_rdata(mshr_16_io_slave_rdata),
    .io_slave_wdata(mshr_16_io_slave_wdata),
    .io_master_req_valid(mshr_16_io_master_req_valid),
    .io_master_req_ready(mshr_16_io_master_req_ready),
    .io_master_req_is_write(mshr_16_io_master_req_is_write),
    .io_master_req_addr(mshr_16_io_master_req_addr),
    .io_master_req_mask(mshr_16_io_master_req_mask),
    .io_master_req_data(mshr_16_io_master_req_data),
    .io_master_resp_valid(mshr_16_io_master_resp_valid),
    .io_master_resp_bits(mshr_16_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_17 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_17_clock),
    .reset(mshr_17_reset),
    .io_enable(mshr_17_io_enable),
    .io_slave_wen(mshr_17_io_slave_wen),
    .io_slave_addr(mshr_17_io_slave_addr),
    .io_slave_rdata(mshr_17_io_slave_rdata),
    .io_slave_wdata(mshr_17_io_slave_wdata),
    .io_master_req_valid(mshr_17_io_master_req_valid),
    .io_master_req_ready(mshr_17_io_master_req_ready),
    .io_master_req_is_write(mshr_17_io_master_req_is_write),
    .io_master_req_addr(mshr_17_io_master_req_addr),
    .io_master_req_mask(mshr_17_io_master_req_mask),
    .io_master_req_data(mshr_17_io_master_req_data),
    .io_master_resp_valid(mshr_17_io_master_resp_valid),
    .io_master_resp_bits(mshr_17_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_18 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_18_clock),
    .reset(mshr_18_reset),
    .io_enable(mshr_18_io_enable),
    .io_slave_wen(mshr_18_io_slave_wen),
    .io_slave_addr(mshr_18_io_slave_addr),
    .io_slave_rdata(mshr_18_io_slave_rdata),
    .io_slave_wdata(mshr_18_io_slave_wdata),
    .io_master_req_valid(mshr_18_io_master_req_valid),
    .io_master_req_ready(mshr_18_io_master_req_ready),
    .io_master_req_is_write(mshr_18_io_master_req_is_write),
    .io_master_req_addr(mshr_18_io_master_req_addr),
    .io_master_req_mask(mshr_18_io_master_req_mask),
    .io_master_req_data(mshr_18_io_master_req_data),
    .io_master_resp_valid(mshr_18_io_master_resp_valid),
    .io_master_resp_bits(mshr_18_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_19 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_19_clock),
    .reset(mshr_19_reset),
    .io_enable(mshr_19_io_enable),
    .io_slave_wen(mshr_19_io_slave_wen),
    .io_slave_addr(mshr_19_io_slave_addr),
    .io_slave_rdata(mshr_19_io_slave_rdata),
    .io_slave_wdata(mshr_19_io_slave_wdata),
    .io_master_req_valid(mshr_19_io_master_req_valid),
    .io_master_req_ready(mshr_19_io_master_req_ready),
    .io_master_req_is_write(mshr_19_io_master_req_is_write),
    .io_master_req_addr(mshr_19_io_master_req_addr),
    .io_master_req_mask(mshr_19_io_master_req_mask),
    .io_master_req_data(mshr_19_io_master_req_data),
    .io_master_resp_valid(mshr_19_io_master_resp_valid),
    .io_master_resp_bits(mshr_19_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_20 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_20_clock),
    .reset(mshr_20_reset),
    .io_enable(mshr_20_io_enable),
    .io_slave_wen(mshr_20_io_slave_wen),
    .io_slave_addr(mshr_20_io_slave_addr),
    .io_slave_rdata(mshr_20_io_slave_rdata),
    .io_slave_wdata(mshr_20_io_slave_wdata),
    .io_master_req_valid(mshr_20_io_master_req_valid),
    .io_master_req_ready(mshr_20_io_master_req_ready),
    .io_master_req_is_write(mshr_20_io_master_req_is_write),
    .io_master_req_addr(mshr_20_io_master_req_addr),
    .io_master_req_mask(mshr_20_io_master_req_mask),
    .io_master_req_data(mshr_20_io_master_req_data),
    .io_master_resp_valid(mshr_20_io_master_resp_valid),
    .io_master_resp_bits(mshr_20_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_21 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_21_clock),
    .reset(mshr_21_reset),
    .io_enable(mshr_21_io_enable),
    .io_slave_wen(mshr_21_io_slave_wen),
    .io_slave_addr(mshr_21_io_slave_addr),
    .io_slave_rdata(mshr_21_io_slave_rdata),
    .io_slave_wdata(mshr_21_io_slave_wdata),
    .io_master_req_valid(mshr_21_io_master_req_valid),
    .io_master_req_ready(mshr_21_io_master_req_ready),
    .io_master_req_is_write(mshr_21_io_master_req_is_write),
    .io_master_req_addr(mshr_21_io_master_req_addr),
    .io_master_req_mask(mshr_21_io_master_req_mask),
    .io_master_req_data(mshr_21_io_master_req_data),
    .io_master_resp_valid(mshr_21_io_master_resp_valid),
    .io_master_resp_bits(mshr_21_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_22 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_22_clock),
    .reset(mshr_22_reset),
    .io_enable(mshr_22_io_enable),
    .io_slave_wen(mshr_22_io_slave_wen),
    .io_slave_addr(mshr_22_io_slave_addr),
    .io_slave_rdata(mshr_22_io_slave_rdata),
    .io_slave_wdata(mshr_22_io_slave_wdata),
    .io_master_req_valid(mshr_22_io_master_req_valid),
    .io_master_req_ready(mshr_22_io_master_req_ready),
    .io_master_req_is_write(mshr_22_io_master_req_is_write),
    .io_master_req_addr(mshr_22_io_master_req_addr),
    .io_master_req_mask(mshr_22_io_master_req_mask),
    .io_master_req_data(mshr_22_io_master_req_data),
    .io_master_resp_valid(mshr_22_io_master_resp_valid),
    .io_master_resp_bits(mshr_22_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_23 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_23_clock),
    .reset(mshr_23_reset),
    .io_enable(mshr_23_io_enable),
    .io_slave_wen(mshr_23_io_slave_wen),
    .io_slave_addr(mshr_23_io_slave_addr),
    .io_slave_rdata(mshr_23_io_slave_rdata),
    .io_slave_wdata(mshr_23_io_slave_wdata),
    .io_master_req_valid(mshr_23_io_master_req_valid),
    .io_master_req_ready(mshr_23_io_master_req_ready),
    .io_master_req_is_write(mshr_23_io_master_req_is_write),
    .io_master_req_addr(mshr_23_io_master_req_addr),
    .io_master_req_mask(mshr_23_io_master_req_mask),
    .io_master_req_data(mshr_23_io_master_req_data),
    .io_master_resp_valid(mshr_23_io_master_resp_valid),
    .io_master_resp_bits(mshr_23_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_24 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_24_clock),
    .reset(mshr_24_reset),
    .io_enable(mshr_24_io_enable),
    .io_slave_wen(mshr_24_io_slave_wen),
    .io_slave_addr(mshr_24_io_slave_addr),
    .io_slave_rdata(mshr_24_io_slave_rdata),
    .io_slave_wdata(mshr_24_io_slave_wdata),
    .io_master_req_valid(mshr_24_io_master_req_valid),
    .io_master_req_ready(mshr_24_io_master_req_ready),
    .io_master_req_is_write(mshr_24_io_master_req_is_write),
    .io_master_req_addr(mshr_24_io_master_req_addr),
    .io_master_req_mask(mshr_24_io_master_req_mask),
    .io_master_req_data(mshr_24_io_master_req_data),
    .io_master_resp_valid(mshr_24_io_master_resp_valid),
    .io_master_resp_bits(mshr_24_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_25 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_25_clock),
    .reset(mshr_25_reset),
    .io_enable(mshr_25_io_enable),
    .io_slave_wen(mshr_25_io_slave_wen),
    .io_slave_addr(mshr_25_io_slave_addr),
    .io_slave_rdata(mshr_25_io_slave_rdata),
    .io_slave_wdata(mshr_25_io_slave_wdata),
    .io_master_req_valid(mshr_25_io_master_req_valid),
    .io_master_req_ready(mshr_25_io_master_req_ready),
    .io_master_req_is_write(mshr_25_io_master_req_is_write),
    .io_master_req_addr(mshr_25_io_master_req_addr),
    .io_master_req_mask(mshr_25_io_master_req_mask),
    .io_master_req_data(mshr_25_io_master_req_data),
    .io_master_resp_valid(mshr_25_io_master_resp_valid),
    .io_master_resp_bits(mshr_25_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_26 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_26_clock),
    .reset(mshr_26_reset),
    .io_enable(mshr_26_io_enable),
    .io_slave_wen(mshr_26_io_slave_wen),
    .io_slave_addr(mshr_26_io_slave_addr),
    .io_slave_rdata(mshr_26_io_slave_rdata),
    .io_slave_wdata(mshr_26_io_slave_wdata),
    .io_master_req_valid(mshr_26_io_master_req_valid),
    .io_master_req_ready(mshr_26_io_master_req_ready),
    .io_master_req_is_write(mshr_26_io_master_req_is_write),
    .io_master_req_addr(mshr_26_io_master_req_addr),
    .io_master_req_mask(mshr_26_io_master_req_mask),
    .io_master_req_data(mshr_26_io_master_req_data),
    .io_master_resp_valid(mshr_26_io_master_resp_valid),
    .io_master_resp_bits(mshr_26_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_27 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_27_clock),
    .reset(mshr_27_reset),
    .io_enable(mshr_27_io_enable),
    .io_slave_wen(mshr_27_io_slave_wen),
    .io_slave_addr(mshr_27_io_slave_addr),
    .io_slave_rdata(mshr_27_io_slave_rdata),
    .io_slave_wdata(mshr_27_io_slave_wdata),
    .io_master_req_valid(mshr_27_io_master_req_valid),
    .io_master_req_ready(mshr_27_io_master_req_ready),
    .io_master_req_is_write(mshr_27_io_master_req_is_write),
    .io_master_req_addr(mshr_27_io_master_req_addr),
    .io_master_req_mask(mshr_27_io_master_req_mask),
    .io_master_req_data(mshr_27_io_master_req_data),
    .io_master_resp_valid(mshr_27_io_master_resp_valid),
    .io_master_resp_bits(mshr_27_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_28 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_28_clock),
    .reset(mshr_28_reset),
    .io_enable(mshr_28_io_enable),
    .io_slave_wen(mshr_28_io_slave_wen),
    .io_slave_addr(mshr_28_io_slave_addr),
    .io_slave_rdata(mshr_28_io_slave_rdata),
    .io_slave_wdata(mshr_28_io_slave_wdata),
    .io_master_req_valid(mshr_28_io_master_req_valid),
    .io_master_req_ready(mshr_28_io_master_req_ready),
    .io_master_req_is_write(mshr_28_io_master_req_is_write),
    .io_master_req_addr(mshr_28_io_master_req_addr),
    .io_master_req_mask(mshr_28_io_master_req_mask),
    .io_master_req_data(mshr_28_io_master_req_data),
    .io_master_resp_valid(mshr_28_io_master_resp_valid),
    .io_master_resp_bits(mshr_28_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_29 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_29_clock),
    .reset(mshr_29_reset),
    .io_enable(mshr_29_io_enable),
    .io_slave_wen(mshr_29_io_slave_wen),
    .io_slave_addr(mshr_29_io_slave_addr),
    .io_slave_rdata(mshr_29_io_slave_rdata),
    .io_slave_wdata(mshr_29_io_slave_wdata),
    .io_master_req_valid(mshr_29_io_master_req_valid),
    .io_master_req_ready(mshr_29_io_master_req_ready),
    .io_master_req_is_write(mshr_29_io_master_req_is_write),
    .io_master_req_addr(mshr_29_io_master_req_addr),
    .io_master_req_mask(mshr_29_io_master_req_mask),
    .io_master_req_data(mshr_29_io_master_req_data),
    .io_master_resp_valid(mshr_29_io_master_resp_valid),
    .io_master_resp_bits(mshr_29_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_30 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_30_clock),
    .reset(mshr_30_reset),
    .io_enable(mshr_30_io_enable),
    .io_slave_wen(mshr_30_io_slave_wen),
    .io_slave_addr(mshr_30_io_slave_addr),
    .io_slave_rdata(mshr_30_io_slave_rdata),
    .io_slave_wdata(mshr_30_io_slave_wdata),
    .io_master_req_valid(mshr_30_io_master_req_valid),
    .io_master_req_ready(mshr_30_io_master_req_ready),
    .io_master_req_is_write(mshr_30_io_master_req_is_write),
    .io_master_req_addr(mshr_30_io_master_req_addr),
    .io_master_req_mask(mshr_30_io_master_req_mask),
    .io_master_req_data(mshr_30_io_master_req_data),
    .io_master_resp_valid(mshr_30_io_master_resp_valid),
    .io_master_resp_bits(mshr_30_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_31 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_31_clock),
    .reset(mshr_31_reset),
    .io_enable(mshr_31_io_enable),
    .io_slave_wen(mshr_31_io_slave_wen),
    .io_slave_addr(mshr_31_io_slave_addr),
    .io_slave_rdata(mshr_31_io_slave_rdata),
    .io_slave_wdata(mshr_31_io_slave_wdata),
    .io_master_req_valid(mshr_31_io_master_req_valid),
    .io_master_req_ready(mshr_31_io_master_req_ready),
    .io_master_req_is_write(mshr_31_io_master_req_is_write),
    .io_master_req_addr(mshr_31_io_master_req_addr),
    .io_master_req_mask(mshr_31_io_master_req_mask),
    .io_master_req_data(mshr_31_io_master_req_data),
    .io_master_resp_valid(mshr_31_io_master_resp_valid),
    .io_master_resp_bits(mshr_31_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_32 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_32_clock),
    .reset(mshr_32_reset),
    .io_enable(mshr_32_io_enable),
    .io_slave_wen(mshr_32_io_slave_wen),
    .io_slave_addr(mshr_32_io_slave_addr),
    .io_slave_rdata(mshr_32_io_slave_rdata),
    .io_slave_wdata(mshr_32_io_slave_wdata),
    .io_master_req_valid(mshr_32_io_master_req_valid),
    .io_master_req_ready(mshr_32_io_master_req_ready),
    .io_master_req_is_write(mshr_32_io_master_req_is_write),
    .io_master_req_addr(mshr_32_io_master_req_addr),
    .io_master_req_mask(mshr_32_io_master_req_mask),
    .io_master_req_data(mshr_32_io_master_req_data),
    .io_master_resp_valid(mshr_32_io_master_resp_valid),
    .io_master_resp_bits(mshr_32_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_33 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_33_clock),
    .reset(mshr_33_reset),
    .io_enable(mshr_33_io_enable),
    .io_slave_wen(mshr_33_io_slave_wen),
    .io_slave_addr(mshr_33_io_slave_addr),
    .io_slave_rdata(mshr_33_io_slave_rdata),
    .io_slave_wdata(mshr_33_io_slave_wdata),
    .io_master_req_valid(mshr_33_io_master_req_valid),
    .io_master_req_ready(mshr_33_io_master_req_ready),
    .io_master_req_is_write(mshr_33_io_master_req_is_write),
    .io_master_req_addr(mshr_33_io_master_req_addr),
    .io_master_req_mask(mshr_33_io_master_req_mask),
    .io_master_req_data(mshr_33_io_master_req_data),
    .io_master_resp_valid(mshr_33_io_master_resp_valid),
    .io_master_resp_bits(mshr_33_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_34 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_34_clock),
    .reset(mshr_34_reset),
    .io_enable(mshr_34_io_enable),
    .io_slave_wen(mshr_34_io_slave_wen),
    .io_slave_addr(mshr_34_io_slave_addr),
    .io_slave_rdata(mshr_34_io_slave_rdata),
    .io_slave_wdata(mshr_34_io_slave_wdata),
    .io_master_req_valid(mshr_34_io_master_req_valid),
    .io_master_req_ready(mshr_34_io_master_req_ready),
    .io_master_req_is_write(mshr_34_io_master_req_is_write),
    .io_master_req_addr(mshr_34_io_master_req_addr),
    .io_master_req_mask(mshr_34_io_master_req_mask),
    .io_master_req_data(mshr_34_io_master_req_data),
    .io_master_resp_valid(mshr_34_io_master_resp_valid),
    .io_master_resp_bits(mshr_34_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_35 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_35_clock),
    .reset(mshr_35_reset),
    .io_enable(mshr_35_io_enable),
    .io_slave_wen(mshr_35_io_slave_wen),
    .io_slave_addr(mshr_35_io_slave_addr),
    .io_slave_rdata(mshr_35_io_slave_rdata),
    .io_slave_wdata(mshr_35_io_slave_wdata),
    .io_master_req_valid(mshr_35_io_master_req_valid),
    .io_master_req_ready(mshr_35_io_master_req_ready),
    .io_master_req_is_write(mshr_35_io_master_req_is_write),
    .io_master_req_addr(mshr_35_io_master_req_addr),
    .io_master_req_mask(mshr_35_io_master_req_mask),
    .io_master_req_data(mshr_35_io_master_req_data),
    .io_master_resp_valid(mshr_35_io_master_resp_valid),
    .io_master_resp_bits(mshr_35_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_36 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_36_clock),
    .reset(mshr_36_reset),
    .io_enable(mshr_36_io_enable),
    .io_slave_wen(mshr_36_io_slave_wen),
    .io_slave_addr(mshr_36_io_slave_addr),
    .io_slave_rdata(mshr_36_io_slave_rdata),
    .io_slave_wdata(mshr_36_io_slave_wdata),
    .io_master_req_valid(mshr_36_io_master_req_valid),
    .io_master_req_ready(mshr_36_io_master_req_ready),
    .io_master_req_is_write(mshr_36_io_master_req_is_write),
    .io_master_req_addr(mshr_36_io_master_req_addr),
    .io_master_req_mask(mshr_36_io_master_req_mask),
    .io_master_req_data(mshr_36_io_master_req_data),
    .io_master_resp_valid(mshr_36_io_master_resp_valid),
    .io_master_resp_bits(mshr_36_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_37 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_37_clock),
    .reset(mshr_37_reset),
    .io_enable(mshr_37_io_enable),
    .io_slave_wen(mshr_37_io_slave_wen),
    .io_slave_addr(mshr_37_io_slave_addr),
    .io_slave_rdata(mshr_37_io_slave_rdata),
    .io_slave_wdata(mshr_37_io_slave_wdata),
    .io_master_req_valid(mshr_37_io_master_req_valid),
    .io_master_req_ready(mshr_37_io_master_req_ready),
    .io_master_req_is_write(mshr_37_io_master_req_is_write),
    .io_master_req_addr(mshr_37_io_master_req_addr),
    .io_master_req_mask(mshr_37_io_master_req_mask),
    .io_master_req_data(mshr_37_io_master_req_data),
    .io_master_resp_valid(mshr_37_io_master_resp_valid),
    .io_master_resp_bits(mshr_37_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_38 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_38_clock),
    .reset(mshr_38_reset),
    .io_enable(mshr_38_io_enable),
    .io_slave_wen(mshr_38_io_slave_wen),
    .io_slave_addr(mshr_38_io_slave_addr),
    .io_slave_rdata(mshr_38_io_slave_rdata),
    .io_slave_wdata(mshr_38_io_slave_wdata),
    .io_master_req_valid(mshr_38_io_master_req_valid),
    .io_master_req_ready(mshr_38_io_master_req_ready),
    .io_master_req_is_write(mshr_38_io_master_req_is_write),
    .io_master_req_addr(mshr_38_io_master_req_addr),
    .io_master_req_mask(mshr_38_io_master_req_mask),
    .io_master_req_data(mshr_38_io_master_req_data),
    .io_master_resp_valid(mshr_38_io_master_resp_valid),
    .io_master_resp_bits(mshr_38_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_39 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_39_clock),
    .reset(mshr_39_reset),
    .io_enable(mshr_39_io_enable),
    .io_slave_wen(mshr_39_io_slave_wen),
    .io_slave_addr(mshr_39_io_slave_addr),
    .io_slave_rdata(mshr_39_io_slave_rdata),
    .io_slave_wdata(mshr_39_io_slave_wdata),
    .io_master_req_valid(mshr_39_io_master_req_valid),
    .io_master_req_ready(mshr_39_io_master_req_ready),
    .io_master_req_is_write(mshr_39_io_master_req_is_write),
    .io_master_req_addr(mshr_39_io_master_req_addr),
    .io_master_req_mask(mshr_39_io_master_req_mask),
    .io_master_req_data(mshr_39_io_master_req_data),
    .io_master_resp_valid(mshr_39_io_master_resp_valid),
    .io_master_resp_bits(mshr_39_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_40 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_40_clock),
    .reset(mshr_40_reset),
    .io_enable(mshr_40_io_enable),
    .io_slave_wen(mshr_40_io_slave_wen),
    .io_slave_addr(mshr_40_io_slave_addr),
    .io_slave_rdata(mshr_40_io_slave_rdata),
    .io_slave_wdata(mshr_40_io_slave_wdata),
    .io_master_req_valid(mshr_40_io_master_req_valid),
    .io_master_req_ready(mshr_40_io_master_req_ready),
    .io_master_req_is_write(mshr_40_io_master_req_is_write),
    .io_master_req_addr(mshr_40_io_master_req_addr),
    .io_master_req_mask(mshr_40_io_master_req_mask),
    .io_master_req_data(mshr_40_io_master_req_data),
    .io_master_resp_valid(mshr_40_io_master_resp_valid),
    .io_master_resp_bits(mshr_40_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_41 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_41_clock),
    .reset(mshr_41_reset),
    .io_enable(mshr_41_io_enable),
    .io_slave_wen(mshr_41_io_slave_wen),
    .io_slave_addr(mshr_41_io_slave_addr),
    .io_slave_rdata(mshr_41_io_slave_rdata),
    .io_slave_wdata(mshr_41_io_slave_wdata),
    .io_master_req_valid(mshr_41_io_master_req_valid),
    .io_master_req_ready(mshr_41_io_master_req_ready),
    .io_master_req_is_write(mshr_41_io_master_req_is_write),
    .io_master_req_addr(mshr_41_io_master_req_addr),
    .io_master_req_mask(mshr_41_io_master_req_mask),
    .io_master_req_data(mshr_41_io_master_req_data),
    .io_master_resp_valid(mshr_41_io_master_resp_valid),
    .io_master_resp_bits(mshr_41_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_42 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_42_clock),
    .reset(mshr_42_reset),
    .io_enable(mshr_42_io_enable),
    .io_slave_wen(mshr_42_io_slave_wen),
    .io_slave_addr(mshr_42_io_slave_addr),
    .io_slave_rdata(mshr_42_io_slave_rdata),
    .io_slave_wdata(mshr_42_io_slave_wdata),
    .io_master_req_valid(mshr_42_io_master_req_valid),
    .io_master_req_ready(mshr_42_io_master_req_ready),
    .io_master_req_is_write(mshr_42_io_master_req_is_write),
    .io_master_req_addr(mshr_42_io_master_req_addr),
    .io_master_req_mask(mshr_42_io_master_req_mask),
    .io_master_req_data(mshr_42_io_master_req_data),
    .io_master_resp_valid(mshr_42_io_master_resp_valid),
    .io_master_resp_bits(mshr_42_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_43 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_43_clock),
    .reset(mshr_43_reset),
    .io_enable(mshr_43_io_enable),
    .io_slave_wen(mshr_43_io_slave_wen),
    .io_slave_addr(mshr_43_io_slave_addr),
    .io_slave_rdata(mshr_43_io_slave_rdata),
    .io_slave_wdata(mshr_43_io_slave_wdata),
    .io_master_req_valid(mshr_43_io_master_req_valid),
    .io_master_req_ready(mshr_43_io_master_req_ready),
    .io_master_req_is_write(mshr_43_io_master_req_is_write),
    .io_master_req_addr(mshr_43_io_master_req_addr),
    .io_master_req_mask(mshr_43_io_master_req_mask),
    .io_master_req_data(mshr_43_io_master_req_data),
    .io_master_resp_valid(mshr_43_io_master_resp_valid),
    .io_master_resp_bits(mshr_43_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_44 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_44_clock),
    .reset(mshr_44_reset),
    .io_enable(mshr_44_io_enable),
    .io_slave_wen(mshr_44_io_slave_wen),
    .io_slave_addr(mshr_44_io_slave_addr),
    .io_slave_rdata(mshr_44_io_slave_rdata),
    .io_slave_wdata(mshr_44_io_slave_wdata),
    .io_master_req_valid(mshr_44_io_master_req_valid),
    .io_master_req_ready(mshr_44_io_master_req_ready),
    .io_master_req_is_write(mshr_44_io_master_req_is_write),
    .io_master_req_addr(mshr_44_io_master_req_addr),
    .io_master_req_mask(mshr_44_io_master_req_mask),
    .io_master_req_data(mshr_44_io_master_req_data),
    .io_master_resp_valid(mshr_44_io_master_resp_valid),
    .io_master_resp_bits(mshr_44_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_45 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_45_clock),
    .reset(mshr_45_reset),
    .io_enable(mshr_45_io_enable),
    .io_slave_wen(mshr_45_io_slave_wen),
    .io_slave_addr(mshr_45_io_slave_addr),
    .io_slave_rdata(mshr_45_io_slave_rdata),
    .io_slave_wdata(mshr_45_io_slave_wdata),
    .io_master_req_valid(mshr_45_io_master_req_valid),
    .io_master_req_ready(mshr_45_io_master_req_ready),
    .io_master_req_is_write(mshr_45_io_master_req_is_write),
    .io_master_req_addr(mshr_45_io_master_req_addr),
    .io_master_req_mask(mshr_45_io_master_req_mask),
    .io_master_req_data(mshr_45_io_master_req_data),
    .io_master_resp_valid(mshr_45_io_master_resp_valid),
    .io_master_resp_bits(mshr_45_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_46 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_46_clock),
    .reset(mshr_46_reset),
    .io_enable(mshr_46_io_enable),
    .io_slave_wen(mshr_46_io_slave_wen),
    .io_slave_addr(mshr_46_io_slave_addr),
    .io_slave_rdata(mshr_46_io_slave_rdata),
    .io_slave_wdata(mshr_46_io_slave_wdata),
    .io_master_req_valid(mshr_46_io_master_req_valid),
    .io_master_req_ready(mshr_46_io_master_req_ready),
    .io_master_req_is_write(mshr_46_io_master_req_is_write),
    .io_master_req_addr(mshr_46_io_master_req_addr),
    .io_master_req_mask(mshr_46_io_master_req_mask),
    .io_master_req_data(mshr_46_io_master_req_data),
    .io_master_resp_valid(mshr_46_io_master_resp_valid),
    .io_master_resp_bits(mshr_46_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_47 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_47_clock),
    .reset(mshr_47_reset),
    .io_enable(mshr_47_io_enable),
    .io_slave_wen(mshr_47_io_slave_wen),
    .io_slave_addr(mshr_47_io_slave_addr),
    .io_slave_rdata(mshr_47_io_slave_rdata),
    .io_slave_wdata(mshr_47_io_slave_wdata),
    .io_master_req_valid(mshr_47_io_master_req_valid),
    .io_master_req_ready(mshr_47_io_master_req_ready),
    .io_master_req_is_write(mshr_47_io_master_req_is_write),
    .io_master_req_addr(mshr_47_io_master_req_addr),
    .io_master_req_mask(mshr_47_io_master_req_mask),
    .io_master_req_data(mshr_47_io_master_req_data),
    .io_master_resp_valid(mshr_47_io_master_resp_valid),
    .io_master_resp_bits(mshr_47_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_48 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_48_clock),
    .reset(mshr_48_reset),
    .io_enable(mshr_48_io_enable),
    .io_slave_wen(mshr_48_io_slave_wen),
    .io_slave_addr(mshr_48_io_slave_addr),
    .io_slave_rdata(mshr_48_io_slave_rdata),
    .io_slave_wdata(mshr_48_io_slave_wdata),
    .io_master_req_valid(mshr_48_io_master_req_valid),
    .io_master_req_ready(mshr_48_io_master_req_ready),
    .io_master_req_is_write(mshr_48_io_master_req_is_write),
    .io_master_req_addr(mshr_48_io_master_req_addr),
    .io_master_req_mask(mshr_48_io_master_req_mask),
    .io_master_req_data(mshr_48_io_master_req_data),
    .io_master_resp_valid(mshr_48_io_master_resp_valid),
    .io_master_resp_bits(mshr_48_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_49 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_49_clock),
    .reset(mshr_49_reset),
    .io_enable(mshr_49_io_enable),
    .io_slave_wen(mshr_49_io_slave_wen),
    .io_slave_addr(mshr_49_io_slave_addr),
    .io_slave_rdata(mshr_49_io_slave_rdata),
    .io_slave_wdata(mshr_49_io_slave_wdata),
    .io_master_req_valid(mshr_49_io_master_req_valid),
    .io_master_req_ready(mshr_49_io_master_req_ready),
    .io_master_req_is_write(mshr_49_io_master_req_is_write),
    .io_master_req_addr(mshr_49_io_master_req_addr),
    .io_master_req_mask(mshr_49_io_master_req_mask),
    .io_master_req_data(mshr_49_io_master_req_data),
    .io_master_resp_valid(mshr_49_io_master_resp_valid),
    .io_master_resp_bits(mshr_49_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_50 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_50_clock),
    .reset(mshr_50_reset),
    .io_enable(mshr_50_io_enable),
    .io_slave_wen(mshr_50_io_slave_wen),
    .io_slave_addr(mshr_50_io_slave_addr),
    .io_slave_rdata(mshr_50_io_slave_rdata),
    .io_slave_wdata(mshr_50_io_slave_wdata),
    .io_master_req_valid(mshr_50_io_master_req_valid),
    .io_master_req_ready(mshr_50_io_master_req_ready),
    .io_master_req_is_write(mshr_50_io_master_req_is_write),
    .io_master_req_addr(mshr_50_io_master_req_addr),
    .io_master_req_mask(mshr_50_io_master_req_mask),
    .io_master_req_data(mshr_50_io_master_req_data),
    .io_master_resp_valid(mshr_50_io_master_resp_valid),
    .io_master_resp_bits(mshr_50_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_51 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_51_clock),
    .reset(mshr_51_reset),
    .io_enable(mshr_51_io_enable),
    .io_slave_wen(mshr_51_io_slave_wen),
    .io_slave_addr(mshr_51_io_slave_addr),
    .io_slave_rdata(mshr_51_io_slave_rdata),
    .io_slave_wdata(mshr_51_io_slave_wdata),
    .io_master_req_valid(mshr_51_io_master_req_valid),
    .io_master_req_ready(mshr_51_io_master_req_ready),
    .io_master_req_is_write(mshr_51_io_master_req_is_write),
    .io_master_req_addr(mshr_51_io_master_req_addr),
    .io_master_req_mask(mshr_51_io_master_req_mask),
    .io_master_req_data(mshr_51_io_master_req_data),
    .io_master_resp_valid(mshr_51_io_master_resp_valid),
    .io_master_resp_bits(mshr_51_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_52 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_52_clock),
    .reset(mshr_52_reset),
    .io_enable(mshr_52_io_enable),
    .io_slave_wen(mshr_52_io_slave_wen),
    .io_slave_addr(mshr_52_io_slave_addr),
    .io_slave_rdata(mshr_52_io_slave_rdata),
    .io_slave_wdata(mshr_52_io_slave_wdata),
    .io_master_req_valid(mshr_52_io_master_req_valid),
    .io_master_req_ready(mshr_52_io_master_req_ready),
    .io_master_req_is_write(mshr_52_io_master_req_is_write),
    .io_master_req_addr(mshr_52_io_master_req_addr),
    .io_master_req_mask(mshr_52_io_master_req_mask),
    .io_master_req_data(mshr_52_io_master_req_data),
    .io_master_resp_valid(mshr_52_io_master_resp_valid),
    .io_master_resp_bits(mshr_52_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_53 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_53_clock),
    .reset(mshr_53_reset),
    .io_enable(mshr_53_io_enable),
    .io_slave_wen(mshr_53_io_slave_wen),
    .io_slave_addr(mshr_53_io_slave_addr),
    .io_slave_rdata(mshr_53_io_slave_rdata),
    .io_slave_wdata(mshr_53_io_slave_wdata),
    .io_master_req_valid(mshr_53_io_master_req_valid),
    .io_master_req_ready(mshr_53_io_master_req_ready),
    .io_master_req_is_write(mshr_53_io_master_req_is_write),
    .io_master_req_addr(mshr_53_io_master_req_addr),
    .io_master_req_mask(mshr_53_io_master_req_mask),
    .io_master_req_data(mshr_53_io_master_req_data),
    .io_master_resp_valid(mshr_53_io_master_resp_valid),
    .io_master_resp_bits(mshr_53_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_54 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_54_clock),
    .reset(mshr_54_reset),
    .io_enable(mshr_54_io_enable),
    .io_slave_wen(mshr_54_io_slave_wen),
    .io_slave_addr(mshr_54_io_slave_addr),
    .io_slave_rdata(mshr_54_io_slave_rdata),
    .io_slave_wdata(mshr_54_io_slave_wdata),
    .io_master_req_valid(mshr_54_io_master_req_valid),
    .io_master_req_ready(mshr_54_io_master_req_ready),
    .io_master_req_is_write(mshr_54_io_master_req_is_write),
    .io_master_req_addr(mshr_54_io_master_req_addr),
    .io_master_req_mask(mshr_54_io_master_req_mask),
    .io_master_req_data(mshr_54_io_master_req_data),
    .io_master_resp_valid(mshr_54_io_master_resp_valid),
    .io_master_resp_bits(mshr_54_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_55 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_55_clock),
    .reset(mshr_55_reset),
    .io_enable(mshr_55_io_enable),
    .io_slave_wen(mshr_55_io_slave_wen),
    .io_slave_addr(mshr_55_io_slave_addr),
    .io_slave_rdata(mshr_55_io_slave_rdata),
    .io_slave_wdata(mshr_55_io_slave_wdata),
    .io_master_req_valid(mshr_55_io_master_req_valid),
    .io_master_req_ready(mshr_55_io_master_req_ready),
    .io_master_req_is_write(mshr_55_io_master_req_is_write),
    .io_master_req_addr(mshr_55_io_master_req_addr),
    .io_master_req_mask(mshr_55_io_master_req_mask),
    .io_master_req_data(mshr_55_io_master_req_data),
    .io_master_resp_valid(mshr_55_io_master_resp_valid),
    .io_master_resp_bits(mshr_55_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_56 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_56_clock),
    .reset(mshr_56_reset),
    .io_enable(mshr_56_io_enable),
    .io_slave_wen(mshr_56_io_slave_wen),
    .io_slave_addr(mshr_56_io_slave_addr),
    .io_slave_rdata(mshr_56_io_slave_rdata),
    .io_slave_wdata(mshr_56_io_slave_wdata),
    .io_master_req_valid(mshr_56_io_master_req_valid),
    .io_master_req_ready(mshr_56_io_master_req_ready),
    .io_master_req_is_write(mshr_56_io_master_req_is_write),
    .io_master_req_addr(mshr_56_io_master_req_addr),
    .io_master_req_mask(mshr_56_io_master_req_mask),
    .io_master_req_data(mshr_56_io_master_req_data),
    .io_master_resp_valid(mshr_56_io_master_resp_valid),
    .io_master_resp_bits(mshr_56_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_57 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_57_clock),
    .reset(mshr_57_reset),
    .io_enable(mshr_57_io_enable),
    .io_slave_wen(mshr_57_io_slave_wen),
    .io_slave_addr(mshr_57_io_slave_addr),
    .io_slave_rdata(mshr_57_io_slave_rdata),
    .io_slave_wdata(mshr_57_io_slave_wdata),
    .io_master_req_valid(mshr_57_io_master_req_valid),
    .io_master_req_ready(mshr_57_io_master_req_ready),
    .io_master_req_is_write(mshr_57_io_master_req_is_write),
    .io_master_req_addr(mshr_57_io_master_req_addr),
    .io_master_req_mask(mshr_57_io_master_req_mask),
    .io_master_req_data(mshr_57_io_master_req_data),
    .io_master_resp_valid(mshr_57_io_master_resp_valid),
    .io_master_resp_bits(mshr_57_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_58 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_58_clock),
    .reset(mshr_58_reset),
    .io_enable(mshr_58_io_enable),
    .io_slave_wen(mshr_58_io_slave_wen),
    .io_slave_addr(mshr_58_io_slave_addr),
    .io_slave_rdata(mshr_58_io_slave_rdata),
    .io_slave_wdata(mshr_58_io_slave_wdata),
    .io_master_req_valid(mshr_58_io_master_req_valid),
    .io_master_req_ready(mshr_58_io_master_req_ready),
    .io_master_req_is_write(mshr_58_io_master_req_is_write),
    .io_master_req_addr(mshr_58_io_master_req_addr),
    .io_master_req_mask(mshr_58_io_master_req_mask),
    .io_master_req_data(mshr_58_io_master_req_data),
    .io_master_resp_valid(mshr_58_io_master_resp_valid),
    .io_master_resp_bits(mshr_58_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_59 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_59_clock),
    .reset(mshr_59_reset),
    .io_enable(mshr_59_io_enable),
    .io_slave_wen(mshr_59_io_slave_wen),
    .io_slave_addr(mshr_59_io_slave_addr),
    .io_slave_rdata(mshr_59_io_slave_rdata),
    .io_slave_wdata(mshr_59_io_slave_wdata),
    .io_master_req_valid(mshr_59_io_master_req_valid),
    .io_master_req_ready(mshr_59_io_master_req_ready),
    .io_master_req_is_write(mshr_59_io_master_req_is_write),
    .io_master_req_addr(mshr_59_io_master_req_addr),
    .io_master_req_mask(mshr_59_io_master_req_mask),
    .io_master_req_data(mshr_59_io_master_req_data),
    .io_master_resp_valid(mshr_59_io_master_resp_valid),
    .io_master_resp_bits(mshr_59_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_60 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_60_clock),
    .reset(mshr_60_reset),
    .io_enable(mshr_60_io_enable),
    .io_slave_wen(mshr_60_io_slave_wen),
    .io_slave_addr(mshr_60_io_slave_addr),
    .io_slave_rdata(mshr_60_io_slave_rdata),
    .io_slave_wdata(mshr_60_io_slave_wdata),
    .io_master_req_valid(mshr_60_io_master_req_valid),
    .io_master_req_ready(mshr_60_io_master_req_ready),
    .io_master_req_is_write(mshr_60_io_master_req_is_write),
    .io_master_req_addr(mshr_60_io_master_req_addr),
    .io_master_req_mask(mshr_60_io_master_req_mask),
    .io_master_req_data(mshr_60_io_master_req_data),
    .io_master_resp_valid(mshr_60_io_master_resp_valid),
    .io_master_resp_bits(mshr_60_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_61 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_61_clock),
    .reset(mshr_61_reset),
    .io_enable(mshr_61_io_enable),
    .io_slave_wen(mshr_61_io_slave_wen),
    .io_slave_addr(mshr_61_io_slave_addr),
    .io_slave_rdata(mshr_61_io_slave_rdata),
    .io_slave_wdata(mshr_61_io_slave_wdata),
    .io_master_req_valid(mshr_61_io_master_req_valid),
    .io_master_req_ready(mshr_61_io_master_req_ready),
    .io_master_req_is_write(mshr_61_io_master_req_is_write),
    .io_master_req_addr(mshr_61_io_master_req_addr),
    .io_master_req_mask(mshr_61_io_master_req_mask),
    .io_master_req_data(mshr_61_io_master_req_data),
    .io_master_resp_valid(mshr_61_io_master_resp_valid),
    .io_master_resp_bits(mshr_61_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_62 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_62_clock),
    .reset(mshr_62_reset),
    .io_enable(mshr_62_io_enable),
    .io_slave_wen(mshr_62_io_slave_wen),
    .io_slave_addr(mshr_62_io_slave_addr),
    .io_slave_rdata(mshr_62_io_slave_rdata),
    .io_slave_wdata(mshr_62_io_slave_wdata),
    .io_master_req_valid(mshr_62_io_master_req_valid),
    .io_master_req_ready(mshr_62_io_master_req_ready),
    .io_master_req_is_write(mshr_62_io_master_req_is_write),
    .io_master_req_addr(mshr_62_io_master_req_addr),
    .io_master_req_mask(mshr_62_io_master_req_mask),
    .io_master_req_data(mshr_62_io_master_req_data),
    .io_master_resp_valid(mshr_62_io_master_resp_valid),
    .io_master_resp_bits(mshr_62_io_master_resp_bits)
  );
  DMAFakeMSHR mshr_63 ( // @[AXI4FakeDMA.scala 149:44]
    .clock(mshr_63_clock),
    .reset(mshr_63_reset),
    .io_enable(mshr_63_io_enable),
    .io_slave_wen(mshr_63_io_slave_wen),
    .io_slave_addr(mshr_63_io_slave_addr),
    .io_slave_rdata(mshr_63_io_slave_rdata),
    .io_slave_wdata(mshr_63_io_slave_wdata),
    .io_master_req_valid(mshr_63_io_master_req_valid),
    .io_master_req_ready(mshr_63_io_master_req_ready),
    .io_master_req_is_write(mshr_63_io_master_req_is_write),
    .io_master_req_addr(mshr_63_io_master_req_addr),
    .io_master_req_mask(mshr_63_io_master_req_mask),
    .io_master_req_data(mshr_63_io_master_req_data),
    .io_master_resp_valid(mshr_63_io_master_resp_valid),
    .io_master_resp_bits(mshr_63_io_master_resp_bits)
  );
  assign auto_dma_out_awvalid = w_valid ? 1'h0 : |_bundleOut_0_awvalid_T; // @[AXI4FakeDMA.scala 199:18 222:20 223:20]
  assign auto_dma_out_awid = {{2'd0}, _bundleOut_0_awid_T_16}; // @[Nodes.scala 1207:84 AXI4FakeDMA.scala 201:20]
  assign auto_dma_out_awaddr = out_write_req_addr[37:0]; // @[Nodes.scala 1207:84 AXI4FakeDMA.scala 202:22]
  assign auto_dma_out_wvalid = w_valid; // @[Nodes.scala 1207:84 AXI4FakeDMA.scala 228:17]
  assign auto_dma_out_wdata = beatCount ? w_data[511:256] : w_data[255:0]; // @[AXI4FakeDMA.scala 230:{21,21}]
  assign auto_dma_out_wstrb = beatCount ? w_mask[63:32] : w_mask[31:0]; // @[AXI4FakeDMA.scala 231:{21,21}]
  assign auto_dma_out_wlast = beatCount; // @[AXI4FakeDMA.scala 232:34]
  assign auto_dma_out_arvalid = |_bundleOut_0_arvalid_T; // @[AXI4FakeDMA.scala 187:41]
  assign auto_dma_out_arid = {{2'd0}, _bundleOut_0_arid_T_16}; // @[Nodes.scala 1207:84 AXI4FakeDMA.scala 189:20]
  assign auto_dma_out_araddr = out_read_req_addr[37:0]; // @[Nodes.scala 1207:84 AXI4FakeDMA.scala 190:22]
  assign auto_in_awready = in_awready; // @[LazyModule.scala 309:16]
  assign auto_in_wready = in_wready; // @[LazyModule.scala 309:16]
  assign auto_in_bvalid = in_bvalid; // @[LazyModule.scala 309:16]
  assign auto_in_bid = in_bid; // @[LazyModule.scala 309:16]
  assign auto_in_bresp = in_bresp; // @[LazyModule.scala 309:16]
  assign auto_in_arready = in_arready; // @[LazyModule.scala 309:16]
  assign auto_in_rvalid = in_rvalid; // @[LazyModule.scala 309:16]
  assign auto_in_rid = in_rid; // @[LazyModule.scala 309:16]
  assign auto_in_rdata = in_rdata; // @[LazyModule.scala 309:16]
  assign auto_in_rresp = in_bresp; // @[LazyModule.scala 309:16]
  assign auto_in_rlast = in_rlast; // @[LazyModule.scala 309:16]
  assign mshr_0_clock = clock;
  assign mshr_0_reset = reset;
  assign mshr_0_io_enable = enable[0]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_0_io_slave_wen = _T_2 & reqWriteIdx == 7'h0 & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_0_io_slave_addr = _T_2 & reqWriteIdx == 7'h0 & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_0_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_0_io_master_req_ready = read_fire | write_fire; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_0_io_master_resp_valid = read_resp_fire | write_resp_fire; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_0_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_1_clock = clock;
  assign mshr_1_reset = reset;
  assign mshr_1_io_enable = enable[1]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_1_io_slave_wen = _T_2 & reqWriteIdx == 7'h1 & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_1_io_slave_addr = _T_2 & reqWriteIdx == 7'h1 & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_1_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_1_io_master_req_ready = read_fire_1 | write_fire_1; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_1_io_master_resp_valid = read_resp_fire_1 | write_resp_fire_1; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_1_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_2_clock = clock;
  assign mshr_2_reset = reset;
  assign mshr_2_io_enable = enable[2]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_2_io_slave_wen = _T_2 & reqWriteIdx == 7'h2 & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_2_io_slave_addr = _T_2 & reqWriteIdx == 7'h2 & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_2_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_2_io_master_req_ready = read_fire_2 | write_fire_2; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_2_io_master_resp_valid = read_resp_fire_2 | write_resp_fire_2; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_2_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_3_clock = clock;
  assign mshr_3_reset = reset;
  assign mshr_3_io_enable = enable[3]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_3_io_slave_wen = _T_2 & reqWriteIdx == 7'h3 & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_3_io_slave_addr = _T_2 & reqWriteIdx == 7'h3 & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_3_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_3_io_master_req_ready = read_fire_3 | write_fire_3; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_3_io_master_resp_valid = read_resp_fire_3 | write_resp_fire_3; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_3_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_4_clock = clock;
  assign mshr_4_reset = reset;
  assign mshr_4_io_enable = enable[4]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_4_io_slave_wen = _T_2 & reqWriteIdx == 7'h4 & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_4_io_slave_addr = _T_2 & reqWriteIdx == 7'h4 & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_4_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_4_io_master_req_ready = read_fire_4 | write_fire_4; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_4_io_master_resp_valid = read_resp_fire_4 | write_resp_fire_4; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_4_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_5_clock = clock;
  assign mshr_5_reset = reset;
  assign mshr_5_io_enable = enable[5]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_5_io_slave_wen = _T_2 & reqWriteIdx == 7'h5 & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_5_io_slave_addr = _T_2 & reqWriteIdx == 7'h5 & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_5_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_5_io_master_req_ready = read_fire_5 | write_fire_5; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_5_io_master_resp_valid = read_resp_fire_5 | write_resp_fire_5; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_5_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_6_clock = clock;
  assign mshr_6_reset = reset;
  assign mshr_6_io_enable = enable[6]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_6_io_slave_wen = _T_2 & reqWriteIdx == 7'h6 & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_6_io_slave_addr = _T_2 & reqWriteIdx == 7'h6 & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_6_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_6_io_master_req_ready = read_fire_6 | write_fire_6; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_6_io_master_resp_valid = read_resp_fire_6 | write_resp_fire_6; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_6_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_7_clock = clock;
  assign mshr_7_reset = reset;
  assign mshr_7_io_enable = enable[7]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_7_io_slave_wen = _T_2 & reqWriteIdx == 7'h7 & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_7_io_slave_addr = _T_2 & reqWriteIdx == 7'h7 & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_7_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_7_io_master_req_ready = read_fire_7 | write_fire_7; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_7_io_master_resp_valid = read_resp_fire_7 | write_resp_fire_7; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_7_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_8_clock = clock;
  assign mshr_8_reset = reset;
  assign mshr_8_io_enable = enable[8]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_8_io_slave_wen = _T_2 & reqWriteIdx == 7'h8 & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_8_io_slave_addr = _T_2 & reqWriteIdx == 7'h8 & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_8_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_8_io_master_req_ready = read_fire_8 | write_fire_8; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_8_io_master_resp_valid = read_resp_fire_8 | write_resp_fire_8; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_8_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_9_clock = clock;
  assign mshr_9_reset = reset;
  assign mshr_9_io_enable = enable[9]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_9_io_slave_wen = _T_2 & reqWriteIdx == 7'h9 & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_9_io_slave_addr = _T_2 & reqWriteIdx == 7'h9 & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_9_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_9_io_master_req_ready = read_fire_9 | write_fire_9; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_9_io_master_resp_valid = read_resp_fire_9 | write_resp_fire_9; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_9_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_10_clock = clock;
  assign mshr_10_reset = reset;
  assign mshr_10_io_enable = enable[10]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_10_io_slave_wen = _T_2 & reqWriteIdx == 7'ha & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_10_io_slave_addr = _T_2 & reqWriteIdx == 7'ha & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_10_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_10_io_master_req_ready = read_fire_10 | write_fire_10; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_10_io_master_resp_valid = read_resp_fire_10 | write_resp_fire_10; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_10_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_11_clock = clock;
  assign mshr_11_reset = reset;
  assign mshr_11_io_enable = enable[11]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_11_io_slave_wen = _T_2 & reqWriteIdx == 7'hb & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_11_io_slave_addr = _T_2 & reqWriteIdx == 7'hb & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_11_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_11_io_master_req_ready = read_fire_11 | write_fire_11; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_11_io_master_resp_valid = read_resp_fire_11 | write_resp_fire_11; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_11_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_12_clock = clock;
  assign mshr_12_reset = reset;
  assign mshr_12_io_enable = enable[12]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_12_io_slave_wen = _T_2 & reqWriteIdx == 7'hc & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_12_io_slave_addr = _T_2 & reqWriteIdx == 7'hc & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_12_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_12_io_master_req_ready = read_fire_12 | write_fire_12; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_12_io_master_resp_valid = read_resp_fire_12 | write_resp_fire_12; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_12_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_13_clock = clock;
  assign mshr_13_reset = reset;
  assign mshr_13_io_enable = enable[13]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_13_io_slave_wen = _T_2 & reqWriteIdx == 7'hd & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_13_io_slave_addr = _T_2 & reqWriteIdx == 7'hd & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_13_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_13_io_master_req_ready = read_fire_13 | write_fire_13; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_13_io_master_resp_valid = read_resp_fire_13 | write_resp_fire_13; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_13_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_14_clock = clock;
  assign mshr_14_reset = reset;
  assign mshr_14_io_enable = enable[14]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_14_io_slave_wen = _T_2 & reqWriteIdx == 7'he & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_14_io_slave_addr = _T_2 & reqWriteIdx == 7'he & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_14_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_14_io_master_req_ready = read_fire_14 | write_fire_14; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_14_io_master_resp_valid = read_resp_fire_14 | write_resp_fire_14; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_14_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_15_clock = clock;
  assign mshr_15_reset = reset;
  assign mshr_15_io_enable = enable[15]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_15_io_slave_wen = _T_2 & reqWriteIdx == 7'hf & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_15_io_slave_addr = _T_2 & reqWriteIdx == 7'hf & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_15_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_15_io_master_req_ready = read_fire_15 | write_fire_15; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_15_io_master_resp_valid = read_resp_fire_15 | write_resp_fire_15; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_15_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_16_clock = clock;
  assign mshr_16_reset = reset;
  assign mshr_16_io_enable = enable[16]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_16_io_slave_wen = _T_2 & reqWriteIdx == 7'h10 & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_16_io_slave_addr = _T_2 & reqWriteIdx == 7'h10 & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_16_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_16_io_master_req_ready = read_fire_16 | write_fire_16; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_16_io_master_resp_valid = read_resp_fire_16 | write_resp_fire_16; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_16_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_17_clock = clock;
  assign mshr_17_reset = reset;
  assign mshr_17_io_enable = enable[17]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_17_io_slave_wen = _T_2 & reqWriteIdx == 7'h11 & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_17_io_slave_addr = _T_2 & reqWriteIdx == 7'h11 & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_17_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_17_io_master_req_ready = read_fire_17 | write_fire_17; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_17_io_master_resp_valid = read_resp_fire_17 | write_resp_fire_17; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_17_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_18_clock = clock;
  assign mshr_18_reset = reset;
  assign mshr_18_io_enable = enable[18]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_18_io_slave_wen = _T_2 & reqWriteIdx == 7'h12 & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_18_io_slave_addr = _T_2 & reqWriteIdx == 7'h12 & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_18_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_18_io_master_req_ready = read_fire_18 | write_fire_18; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_18_io_master_resp_valid = read_resp_fire_18 | write_resp_fire_18; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_18_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_19_clock = clock;
  assign mshr_19_reset = reset;
  assign mshr_19_io_enable = enable[19]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_19_io_slave_wen = _T_2 & reqWriteIdx == 7'h13 & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_19_io_slave_addr = _T_2 & reqWriteIdx == 7'h13 & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_19_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_19_io_master_req_ready = read_fire_19 | write_fire_19; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_19_io_master_resp_valid = read_resp_fire_19 | write_resp_fire_19; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_19_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_20_clock = clock;
  assign mshr_20_reset = reset;
  assign mshr_20_io_enable = enable[20]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_20_io_slave_wen = _T_2 & reqWriteIdx == 7'h14 & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_20_io_slave_addr = _T_2 & reqWriteIdx == 7'h14 & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_20_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_20_io_master_req_ready = read_fire_20 | write_fire_20; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_20_io_master_resp_valid = read_resp_fire_20 | write_resp_fire_20; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_20_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_21_clock = clock;
  assign mshr_21_reset = reset;
  assign mshr_21_io_enable = enable[21]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_21_io_slave_wen = _T_2 & reqWriteIdx == 7'h15 & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_21_io_slave_addr = _T_2 & reqWriteIdx == 7'h15 & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_21_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_21_io_master_req_ready = read_fire_21 | write_fire_21; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_21_io_master_resp_valid = read_resp_fire_21 | write_resp_fire_21; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_21_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_22_clock = clock;
  assign mshr_22_reset = reset;
  assign mshr_22_io_enable = enable[22]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_22_io_slave_wen = _T_2 & reqWriteIdx == 7'h16 & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_22_io_slave_addr = _T_2 & reqWriteIdx == 7'h16 & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_22_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_22_io_master_req_ready = read_fire_22 | write_fire_22; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_22_io_master_resp_valid = read_resp_fire_22 | write_resp_fire_22; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_22_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_23_clock = clock;
  assign mshr_23_reset = reset;
  assign mshr_23_io_enable = enable[23]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_23_io_slave_wen = _T_2 & reqWriteIdx == 7'h17 & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_23_io_slave_addr = _T_2 & reqWriteIdx == 7'h17 & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_23_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_23_io_master_req_ready = read_fire_23 | write_fire_23; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_23_io_master_resp_valid = read_resp_fire_23 | write_resp_fire_23; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_23_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_24_clock = clock;
  assign mshr_24_reset = reset;
  assign mshr_24_io_enable = enable[24]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_24_io_slave_wen = _T_2 & reqWriteIdx == 7'h18 & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_24_io_slave_addr = _T_2 & reqWriteIdx == 7'h18 & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_24_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_24_io_master_req_ready = read_fire_24 | write_fire_24; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_24_io_master_resp_valid = read_resp_fire_24 | write_resp_fire_24; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_24_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_25_clock = clock;
  assign mshr_25_reset = reset;
  assign mshr_25_io_enable = enable[25]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_25_io_slave_wen = _T_2 & reqWriteIdx == 7'h19 & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_25_io_slave_addr = _T_2 & reqWriteIdx == 7'h19 & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_25_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_25_io_master_req_ready = read_fire_25 | write_fire_25; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_25_io_master_resp_valid = read_resp_fire_25 | write_resp_fire_25; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_25_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_26_clock = clock;
  assign mshr_26_reset = reset;
  assign mshr_26_io_enable = enable[26]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_26_io_slave_wen = _T_2 & reqWriteIdx == 7'h1a & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_26_io_slave_addr = _T_2 & reqWriteIdx == 7'h1a & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_26_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_26_io_master_req_ready = read_fire_26 | write_fire_26; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_26_io_master_resp_valid = read_resp_fire_26 | write_resp_fire_26; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_26_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_27_clock = clock;
  assign mshr_27_reset = reset;
  assign mshr_27_io_enable = enable[27]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_27_io_slave_wen = _T_2 & reqWriteIdx == 7'h1b & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_27_io_slave_addr = _T_2 & reqWriteIdx == 7'h1b & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_27_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_27_io_master_req_ready = read_fire_27 | write_fire_27; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_27_io_master_resp_valid = read_resp_fire_27 | write_resp_fire_27; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_27_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_28_clock = clock;
  assign mshr_28_reset = reset;
  assign mshr_28_io_enable = enable[28]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_28_io_slave_wen = _T_2 & reqWriteIdx == 7'h1c & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_28_io_slave_addr = _T_2 & reqWriteIdx == 7'h1c & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_28_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_28_io_master_req_ready = read_fire_28 | write_fire_28; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_28_io_master_resp_valid = read_resp_fire_28 | write_resp_fire_28; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_28_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_29_clock = clock;
  assign mshr_29_reset = reset;
  assign mshr_29_io_enable = enable[29]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_29_io_slave_wen = _T_2 & reqWriteIdx == 7'h1d & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_29_io_slave_addr = _T_2 & reqWriteIdx == 7'h1d & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_29_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_29_io_master_req_ready = read_fire_29 | write_fire_29; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_29_io_master_resp_valid = read_resp_fire_29 | write_resp_fire_29; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_29_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_30_clock = clock;
  assign mshr_30_reset = reset;
  assign mshr_30_io_enable = enable[30]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_30_io_slave_wen = _T_2 & reqWriteIdx == 7'h1e & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_30_io_slave_addr = _T_2 & reqWriteIdx == 7'h1e & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_30_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_30_io_master_req_ready = read_fire_30 | write_fire_30; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_30_io_master_resp_valid = read_resp_fire_30 | write_resp_fire_30; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_30_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_31_clock = clock;
  assign mshr_31_reset = reset;
  assign mshr_31_io_enable = enable[31]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_31_io_slave_wen = _T_2 & reqWriteIdx == 7'h1f & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_31_io_slave_addr = _T_2 & reqWriteIdx == 7'h1f & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_31_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_31_io_master_req_ready = read_fire_31 | write_fire_31; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_31_io_master_resp_valid = read_resp_fire_31 | write_resp_fire_31; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_31_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_32_clock = clock;
  assign mshr_32_reset = reset;
  assign mshr_32_io_enable = enable[32]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_32_io_slave_wen = _T_2 & reqWriteIdx == 7'h20 & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_32_io_slave_addr = _T_2 & reqWriteIdx == 7'h20 & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_32_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_32_io_master_req_ready = read_fire_32 | write_fire_32; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_32_io_master_resp_valid = read_resp_fire_32 | write_resp_fire_32; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_32_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_33_clock = clock;
  assign mshr_33_reset = reset;
  assign mshr_33_io_enable = enable[33]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_33_io_slave_wen = _T_2 & reqWriteIdx == 7'h21 & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_33_io_slave_addr = _T_2 & reqWriteIdx == 7'h21 & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_33_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_33_io_master_req_ready = read_fire_33 | write_fire_33; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_33_io_master_resp_valid = read_resp_fire_33 | write_resp_fire_33; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_33_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_34_clock = clock;
  assign mshr_34_reset = reset;
  assign mshr_34_io_enable = enable[34]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_34_io_slave_wen = _T_2 & reqWriteIdx == 7'h22 & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_34_io_slave_addr = _T_2 & reqWriteIdx == 7'h22 & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_34_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_34_io_master_req_ready = read_fire_34 | write_fire_34; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_34_io_master_resp_valid = read_resp_fire_34 | write_resp_fire_34; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_34_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_35_clock = clock;
  assign mshr_35_reset = reset;
  assign mshr_35_io_enable = enable[35]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_35_io_slave_wen = _T_2 & reqWriteIdx == 7'h23 & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_35_io_slave_addr = _T_2 & reqWriteIdx == 7'h23 & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_35_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_35_io_master_req_ready = read_fire_35 | write_fire_35; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_35_io_master_resp_valid = read_resp_fire_35 | write_resp_fire_35; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_35_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_36_clock = clock;
  assign mshr_36_reset = reset;
  assign mshr_36_io_enable = enable[36]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_36_io_slave_wen = _T_2 & reqWriteIdx == 7'h24 & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_36_io_slave_addr = _T_2 & reqWriteIdx == 7'h24 & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_36_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_36_io_master_req_ready = read_fire_36 | write_fire_36; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_36_io_master_resp_valid = read_resp_fire_36 | write_resp_fire_36; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_36_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_37_clock = clock;
  assign mshr_37_reset = reset;
  assign mshr_37_io_enable = enable[37]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_37_io_slave_wen = _T_2 & reqWriteIdx == 7'h25 & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_37_io_slave_addr = _T_2 & reqWriteIdx == 7'h25 & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_37_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_37_io_master_req_ready = read_fire_37 | write_fire_37; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_37_io_master_resp_valid = read_resp_fire_37 | write_resp_fire_37; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_37_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_38_clock = clock;
  assign mshr_38_reset = reset;
  assign mshr_38_io_enable = enable[38]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_38_io_slave_wen = _T_2 & reqWriteIdx == 7'h26 & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_38_io_slave_addr = _T_2 & reqWriteIdx == 7'h26 & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_38_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_38_io_master_req_ready = read_fire_38 | write_fire_38; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_38_io_master_resp_valid = read_resp_fire_38 | write_resp_fire_38; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_38_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_39_clock = clock;
  assign mshr_39_reset = reset;
  assign mshr_39_io_enable = enable[39]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_39_io_slave_wen = _T_2 & reqWriteIdx == 7'h27 & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_39_io_slave_addr = _T_2 & reqWriteIdx == 7'h27 & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_39_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_39_io_master_req_ready = read_fire_39 | write_fire_39; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_39_io_master_resp_valid = read_resp_fire_39 | write_resp_fire_39; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_39_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_40_clock = clock;
  assign mshr_40_reset = reset;
  assign mshr_40_io_enable = enable[40]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_40_io_slave_wen = _T_2 & reqWriteIdx == 7'h28 & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_40_io_slave_addr = _T_2 & reqWriteIdx == 7'h28 & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_40_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_40_io_master_req_ready = read_fire_40 | write_fire_40; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_40_io_master_resp_valid = read_resp_fire_40 | write_resp_fire_40; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_40_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_41_clock = clock;
  assign mshr_41_reset = reset;
  assign mshr_41_io_enable = enable[41]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_41_io_slave_wen = _T_2 & reqWriteIdx == 7'h29 & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_41_io_slave_addr = _T_2 & reqWriteIdx == 7'h29 & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_41_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_41_io_master_req_ready = read_fire_41 | write_fire_41; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_41_io_master_resp_valid = read_resp_fire_41 | write_resp_fire_41; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_41_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_42_clock = clock;
  assign mshr_42_reset = reset;
  assign mshr_42_io_enable = enable[42]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_42_io_slave_wen = _T_2 & reqWriteIdx == 7'h2a & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_42_io_slave_addr = _T_2 & reqWriteIdx == 7'h2a & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_42_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_42_io_master_req_ready = read_fire_42 | write_fire_42; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_42_io_master_resp_valid = read_resp_fire_42 | write_resp_fire_42; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_42_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_43_clock = clock;
  assign mshr_43_reset = reset;
  assign mshr_43_io_enable = enable[43]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_43_io_slave_wen = _T_2 & reqWriteIdx == 7'h2b & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_43_io_slave_addr = _T_2 & reqWriteIdx == 7'h2b & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_43_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_43_io_master_req_ready = read_fire_43 | write_fire_43; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_43_io_master_resp_valid = read_resp_fire_43 | write_resp_fire_43; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_43_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_44_clock = clock;
  assign mshr_44_reset = reset;
  assign mshr_44_io_enable = enable[44]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_44_io_slave_wen = _T_2 & reqWriteIdx == 7'h2c & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_44_io_slave_addr = _T_2 & reqWriteIdx == 7'h2c & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_44_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_44_io_master_req_ready = read_fire_44 | write_fire_44; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_44_io_master_resp_valid = read_resp_fire_44 | write_resp_fire_44; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_44_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_45_clock = clock;
  assign mshr_45_reset = reset;
  assign mshr_45_io_enable = enable[45]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_45_io_slave_wen = _T_2 & reqWriteIdx == 7'h2d & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_45_io_slave_addr = _T_2 & reqWriteIdx == 7'h2d & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_45_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_45_io_master_req_ready = read_fire_45 | write_fire_45; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_45_io_master_resp_valid = read_resp_fire_45 | write_resp_fire_45; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_45_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_46_clock = clock;
  assign mshr_46_reset = reset;
  assign mshr_46_io_enable = enable[46]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_46_io_slave_wen = _T_2 & reqWriteIdx == 7'h2e & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_46_io_slave_addr = _T_2 & reqWriteIdx == 7'h2e & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_46_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_46_io_master_req_ready = read_fire_46 | write_fire_46; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_46_io_master_resp_valid = read_resp_fire_46 | write_resp_fire_46; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_46_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_47_clock = clock;
  assign mshr_47_reset = reset;
  assign mshr_47_io_enable = enable[47]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_47_io_slave_wen = _T_2 & reqWriteIdx == 7'h2f & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_47_io_slave_addr = _T_2 & reqWriteIdx == 7'h2f & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_47_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_47_io_master_req_ready = read_fire_47 | write_fire_47; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_47_io_master_resp_valid = read_resp_fire_47 | write_resp_fire_47; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_47_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_48_clock = clock;
  assign mshr_48_reset = reset;
  assign mshr_48_io_enable = enable[48]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_48_io_slave_wen = _T_2 & reqWriteIdx == 7'h30 & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_48_io_slave_addr = _T_2 & reqWriteIdx == 7'h30 & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_48_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_48_io_master_req_ready = read_fire_48 | write_fire_48; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_48_io_master_resp_valid = read_resp_fire_48 | write_resp_fire_48; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_48_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_49_clock = clock;
  assign mshr_49_reset = reset;
  assign mshr_49_io_enable = enable[49]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_49_io_slave_wen = _T_2 & reqWriteIdx == 7'h31 & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_49_io_slave_addr = _T_2 & reqWriteIdx == 7'h31 & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_49_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_49_io_master_req_ready = read_fire_49 | write_fire_49; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_49_io_master_resp_valid = read_resp_fire_49 | write_resp_fire_49; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_49_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_50_clock = clock;
  assign mshr_50_reset = reset;
  assign mshr_50_io_enable = enable[50]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_50_io_slave_wen = _T_2 & reqWriteIdx == 7'h32 & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_50_io_slave_addr = _T_2 & reqWriteIdx == 7'h32 & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_50_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_50_io_master_req_ready = read_fire_50 | write_fire_50; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_50_io_master_resp_valid = read_resp_fire_50 | write_resp_fire_50; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_50_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_51_clock = clock;
  assign mshr_51_reset = reset;
  assign mshr_51_io_enable = enable[51]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_51_io_slave_wen = _T_2 & reqWriteIdx == 7'h33 & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_51_io_slave_addr = _T_2 & reqWriteIdx == 7'h33 & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_51_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_51_io_master_req_ready = read_fire_51 | write_fire_51; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_51_io_master_resp_valid = read_resp_fire_51 | write_resp_fire_51; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_51_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_52_clock = clock;
  assign mshr_52_reset = reset;
  assign mshr_52_io_enable = enable[52]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_52_io_slave_wen = _T_2 & reqWriteIdx == 7'h34 & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_52_io_slave_addr = _T_2 & reqWriteIdx == 7'h34 & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_52_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_52_io_master_req_ready = read_fire_52 | write_fire_52; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_52_io_master_resp_valid = read_resp_fire_52 | write_resp_fire_52; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_52_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_53_clock = clock;
  assign mshr_53_reset = reset;
  assign mshr_53_io_enable = enable[53]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_53_io_slave_wen = _T_2 & reqWriteIdx == 7'h35 & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_53_io_slave_addr = _T_2 & reqWriteIdx == 7'h35 & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_53_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_53_io_master_req_ready = read_fire_53 | write_fire_53; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_53_io_master_resp_valid = read_resp_fire_53 | write_resp_fire_53; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_53_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_54_clock = clock;
  assign mshr_54_reset = reset;
  assign mshr_54_io_enable = enable[54]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_54_io_slave_wen = _T_2 & reqWriteIdx == 7'h36 & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_54_io_slave_addr = _T_2 & reqWriteIdx == 7'h36 & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_54_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_54_io_master_req_ready = read_fire_54 | write_fire_54; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_54_io_master_resp_valid = read_resp_fire_54 | write_resp_fire_54; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_54_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_55_clock = clock;
  assign mshr_55_reset = reset;
  assign mshr_55_io_enable = enable[55]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_55_io_slave_wen = _T_2 & reqWriteIdx == 7'h37 & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_55_io_slave_addr = _T_2 & reqWriteIdx == 7'h37 & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_55_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_55_io_master_req_ready = read_fire_55 | write_fire_55; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_55_io_master_resp_valid = read_resp_fire_55 | write_resp_fire_55; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_55_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_56_clock = clock;
  assign mshr_56_reset = reset;
  assign mshr_56_io_enable = enable[56]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_56_io_slave_wen = _T_2 & reqWriteIdx == 7'h38 & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_56_io_slave_addr = _T_2 & reqWriteIdx == 7'h38 & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_56_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_56_io_master_req_ready = read_fire_56 | write_fire_56; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_56_io_master_resp_valid = read_resp_fire_56 | write_resp_fire_56; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_56_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_57_clock = clock;
  assign mshr_57_reset = reset;
  assign mshr_57_io_enable = enable[57]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_57_io_slave_wen = _T_2 & reqWriteIdx == 7'h39 & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_57_io_slave_addr = _T_2 & reqWriteIdx == 7'h39 & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_57_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_57_io_master_req_ready = read_fire_57 | write_fire_57; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_57_io_master_resp_valid = read_resp_fire_57 | write_resp_fire_57; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_57_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_58_clock = clock;
  assign mshr_58_reset = reset;
  assign mshr_58_io_enable = enable[58]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_58_io_slave_wen = _T_2 & reqWriteIdx == 7'h3a & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_58_io_slave_addr = _T_2 & reqWriteIdx == 7'h3a & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_58_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_58_io_master_req_ready = read_fire_58 | write_fire_58; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_58_io_master_resp_valid = read_resp_fire_58 | write_resp_fire_58; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_58_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_59_clock = clock;
  assign mshr_59_reset = reset;
  assign mshr_59_io_enable = enable[59]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_59_io_slave_wen = _T_2 & reqWriteIdx == 7'h3b & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_59_io_slave_addr = _T_2 & reqWriteIdx == 7'h3b & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_59_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_59_io_master_req_ready = read_fire_59 | write_fire_59; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_59_io_master_resp_valid = read_resp_fire_59 | write_resp_fire_59; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_59_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_60_clock = clock;
  assign mshr_60_reset = reset;
  assign mshr_60_io_enable = enable[60]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_60_io_slave_wen = _T_2 & reqWriteIdx == 7'h3c & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_60_io_slave_addr = _T_2 & reqWriteIdx == 7'h3c & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_60_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_60_io_master_req_ready = read_fire_60 | write_fire_60; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_60_io_master_resp_valid = read_resp_fire_60 | write_resp_fire_60; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_60_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_61_clock = clock;
  assign mshr_61_reset = reset;
  assign mshr_61_io_enable = enable[61]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_61_io_slave_wen = _T_2 & reqWriteIdx == 7'h3d & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_61_io_slave_addr = _T_2 & reqWriteIdx == 7'h3d & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_61_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_61_io_master_req_ready = read_fire_61 | write_fire_61; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_61_io_master_resp_valid = read_resp_fire_61 | write_resp_fire_61; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_61_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_62_clock = clock;
  assign mshr_62_reset = reset;
  assign mshr_62_io_enable = enable[62]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_62_io_slave_wen = _T_2 & reqWriteIdx == 7'h3e & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_62_io_slave_addr = _T_2 & reqWriteIdx == 7'h3e & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_62_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_62_io_master_req_ready = read_fire_62 | write_fire_62; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_62_io_master_resp_valid = read_resp_fire_62 | write_resp_fire_62; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_62_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  assign mshr_63_clock = clock;
  assign mshr_63_reset = reset;
  assign mshr_63_io_enable = enable[63]; // @[AXI4FakeDMA.scala 152:21]
  assign mshr_63_io_slave_wen = _T_2 & reqWriteIdx == 7'h3f & ~_GEN_13[13]; // @[AXI4FakeDMA.scala 165:46]
  assign mshr_63_io_slave_addr = _T_2 & reqWriteIdx == 7'h3f & ~_GEN_13[13] ? reqWriteOffset : reqReadOffset; // @[AXI4FakeDMA.scala 123:19 128:19 165:74]
  assign mshr_63_io_slave_wdata = in_wdata; // @[AXI4FakeDMA.scala 129:20 165:74]
  assign mshr_63_io_master_req_ready = read_fire_63 | write_fire_63; // @[AXI4FakeDMA.scala 211:30]
  assign mshr_63_io_master_resp_valid = read_resp_fire_63 | write_resp_fire_63; // @[AXI4FakeDMA.scala 243:36]
  assign mshr_63_io_master_resp_bits = auto_dma_out_rdata; // @[Nodes.scala 1207:84 LazyModule.scala 311:12]
  always @(posedge clock) begin
    if (reset) begin // @[AXI4SlaveModule.scala 95:22]
      state <= 2'h0; // @[AXI4SlaveModule.scala 95:22]
    end else if (2'h0 == state) begin // @[AXI4SlaveModule.scala 97:16]
      if (_T_1) begin // @[AXI4SlaveModule.scala 102:25]
        state <= 2'h2; // @[AXI4SlaveModule.scala 103:15]
      end else if (_T) begin // @[AXI4SlaveModule.scala 99:25]
        state <= 2'h1; // @[AXI4SlaveModule.scala 100:15]
      end
    end else if (2'h1 == state) begin // @[AXI4SlaveModule.scala 97:16]
      if (_T_4 & in_rlast) begin // @[AXI4SlaveModule.scala 107:42]
        state <= 2'h0; // @[AXI4SlaveModule.scala 108:15]
      end
    end else if (2'h2 == state) begin // @[AXI4SlaveModule.scala 97:16]
      state <= _GEN_3;
    end else begin
      state <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      value <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_4) begin // @[AXI4SlaveModule.scala 135:23]
      if (in_rlast) begin // @[AXI4SlaveModule.scala 137:28]
        value <= 8'h0; // @[AXI4SlaveModule.scala 138:17]
      end else begin
        value <= _value_T_1; // @[Counter.scala 78:15]
      end
    end
    if (_T) begin // @[Reg.scala 17:18]
      hold_data <= in_arlen; // @[Reg.scala 17:22]
    end
    if (_T) begin // @[Reg.scala 17:18]
      raddr_hold_data <= in_araddr; // @[Reg.scala 17:22]
    end
    if (_T_1) begin // @[Reg.scala 17:18]
      waddr_hold_data <= in_awaddr; // @[Reg.scala 17:22]
    end
    if (_T_1) begin // @[Reg.scala 17:18]
      bundleIn_0_bid_r <= in_awid; // @[Reg.scala 17:22]
    end
    if (_T) begin // @[Reg.scala 17:18]
      bundleIn_0_rid_r <= in_arid; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[AXI4FakeDMA.scala 151:25]
      enable <= 64'h0; // @[AXI4FakeDMA.scala 151:25]
    end else if (_T_2 & _GEN_13[13]) begin // @[AXI4FakeDMA.scala 169:48]
      enable <= in_wdata; // @[AXI4FakeDMA.scala 170:14]
    end
    if (reset) begin // @[AXI4FakeDMA.scala 215:26]
      w_valid <= 1'h0; // @[AXI4FakeDMA.scala 215:26]
    end else begin
      w_valid <= _GEN_276;
    end
    if (reset) begin // @[AXI4FakeDMA.scala 225:28]
      beatCount <= 1'h0; // @[AXI4FakeDMA.scala 225:28]
    end else if (_T_495) begin // @[AXI4FakeDMA.scala 233:23]
      beatCount <= beatCount + 1'h1; // @[AXI4FakeDMA.scala 234:17]
    end
    if (_write_fire_T) begin // @[Reg.scala 17:18]
      w_mask <= out_write_req_mask; // @[Reg.scala 17:22]
    end
    if (_write_fire_T) begin // @[Reg.scala 17:18]
      w_data <= out_write_req_data; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  value = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  hold_data = _RAND_2[7:0];
  _RAND_3 = {2{`RANDOM}};
  raddr_hold_data = _RAND_3[36:0];
  _RAND_4 = {2{`RANDOM}};
  waddr_hold_data = _RAND_4[36:0];
  _RAND_5 = {1{`RANDOM}};
  bundleIn_0_bid_r = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  bundleIn_0_rid_r = _RAND_6[0:0];
  _RAND_7 = {2{`RANDOM}};
  enable = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  w_valid = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  beatCount = _RAND_9[0:0];
  _RAND_10 = {2{`RANDOM}};
  w_mask = _RAND_10[63:0];
  _RAND_11 = {16{`RANDOM}};
  w_data = _RAND_11[511:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

