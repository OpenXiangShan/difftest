/***************************************************************************************
* Copyright (c) 2020-2023 Institute of Computing Technology, Chinese Academy of Sciences
* Copyright (c) 2020-2021 Peng Cheng Laboratory
*
* DiffTest is licensed under Mulan PSL v2.
* You can use this software according to the terms and conditions of the Mulan PSL v2.
* You may obtain a copy of Mulan PSL v2 at:
*          http://license.coscl.org.cn/MulanPSL2
*
* THIS SOFTWARE IS PROVIDED ON AN "AS IS" BASIS, WITHOUT WARRANTIES OF ANY KIND,
* EITHER EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO NON-INFRINGEMENT,
* MERCHANTABILITY OR FIT FOR A PARTICULAR PURPOSE.
*
* See the Mulan PSL v2 for more details.
***************************************************************************************/

`include "DifftestMacros.v"
module tb_top();

`ifndef TB_NO_DPIC
import "DPI-C" function void set_bin_file(string bin);
import "DPI-C" function void set_flash_bin(string bin);
import "DPI-C" function void set_gcpt_bin(string bin);
import "DPI-C" function void set_diff_ref_so(string diff_so);
import "DPI-C" function void set_no_diff();
import "DPI-C" function void set_max_instrs(int mc);
import "DPI-C" function void get_ipc(longint cycles);
import "DPI-C" function void simv_init();
`ifndef CONFIG_DIFFTEST_DEFERRED_RESULT
import "DPI-C" function int simv_nstep(int step);
`endif // CONFIG_DIFFTEST_DEFERRED_RESULT
`ifdef PALLADIUM
import "DPI-C" function void difftest_checkpoint_list(string path);
import "DPI-C" function byte difftest_ram_reload();
`endif // PALLADIUM
`endif // TB_NO_DPIC

`ifdef PALLADIUM
  `ifdef SYNTHESIS
  `define WIRE_CLK //clock will be generated by ixclkgen
  `endif // SYNTHESIS
`endif // PALLADIUM

`ifdef WIRE_CLK
wire        clock;
`else
reg         clock;
`endif // WIRE_CLK
reg         reset;
reg  [63:0] difftest_logCtrl_begin;
reg  [63:0] difftest_logCtrl_end;
wire [63:0] difftest_logCtrl_level;
wire        difftest_perfCtrl_clean;
wire        difftest_perfCtrl_dump;
wire        difftest_uart_out_valid;
wire [ 7:0] difftest_uart_out_ch;
wire        difftest_uart_in_valid;
wire [ 7:0] difftest_uart_in_ch;
wire [`CONFIG_DIFFTEST_STEPWIDTH - 1:0] difftest_step;

string bin_file;
string flash_bin_file;
string gcpt_bin_file;
string wave_type;
string diff_ref_so;
string ckpt_list;

reg [63:0] max_instrs;
reg [63:0] max_cycles;
reg ckpt_list_en;
reg xs_rst_en;

initial begin
`ifndef WIRE_CLK
  clock = 0;
`endif // WIRE_CLK
  reset = 1;

`ifdef VCS
  // enable waveform
  if ($test$plusargs("dump-wave")) begin
    $value$plusargs("dump-wave=%s", wave_type);
    if (wave_type == "vpd") begin
      $vcdplusfile("simv.vpd");
      $vcdpluson;
    end
`ifdef CONSIDER_FSDB
    else if (wave_type == "fsdb") begin
      $fsdbDumpfile("simv.fsdb");
      $fsdbDumpvars(0,"+mda");
    end
`endif
    else begin
      $display("unknown wave file format, want [vpd, fsdb] but:%s\n", wave_type);
      $finish();
    end
  end
`endif

  // log begin
  if ($test$plusargs("b")) begin
    $value$plusargs("b=%d", difftest_logCtrl_begin);
  end
  else begin
    difftest_logCtrl_begin = 0;
  end
  // log end
  if ($test$plusargs("e")) begin
    $value$plusargs("e=%d", difftest_logCtrl_end);
  end
  else begin
    difftest_logCtrl_end = 0;
  end
`ifndef TB_NO_DPIC
  // workload: bin file
  if ($test$plusargs("workload")) begin
    $value$plusargs("workload=%s", bin_file);
    set_bin_file(bin_file);
  end
  // boot flash image: bin file
  if ($test$plusargs("flash")) begin
    $value$plusargs("flash=%s", flash_bin_file);
    set_flash_bin(flash_bin_file);
  end
  // override gcpt :bin file
  if ($test$plusargs("gcpt-bin")) begin
    $value$plusargs("gcpt-bin=%s", gcpt_bin_file);
    set_gcpt_bin(gcpt_bin_file);
  end
  // diff-test golden model: nemu-so
  if ($test$plusargs("diff")) begin
    $value$plusargs("diff=%s", diff_ref_so);
    set_diff_ref_so(diff_ref_so);
  end
  // disable diff-test
  if ($test$plusargs("no-diff")) begin
    set_no_diff();
  end
  // set checkpoint run list
  if ($test$plusargs("ckpt-list")) begin
    $value$plusargs("ckpt-list=%s", ckpt_list);
    difftest_checkpoint_list(ckpt_list);
    ckpt_list_en = 1;
  end

`endif // TB_NO_DPIC
  // max cycles to execute, no limit for default
  max_cycles = 0;
  if ($test$plusargs("max-cycles")) begin
    $value$plusargs("max-cycles=%d", max_cycles);
    $display("set max cycles: %d", max_cycles);
  end
  // set checkpoint const
  if ($test$plusargs("max-instrs")) begin
    $value$plusargs("max-instrs=%d", max_instrs);
    set_max_instrs(max_instrs);
  end
  else begin
    max_instrs = 0;
  end
end

// Note: reset delay #100 should be larger than RANDOMIZE_DELAY
`ifndef PALLADIUM
initial begin
  #100 reset = 0;
end
`else
reg [7:0] reset_counter;
initial reset_counter = 0;
always @(posedge clock) begin
  if (xs_rst_en) begin
    reset_counter <= 8'd0;
    reset         <= 1'b1;
    $display("soft rst CPU core");
  end 
  else begin
    if (reset && (reset_counter == 8'd100)) begin
      reset <= 1'b0;
      $display("rst unlock");
    end else if (reset) begin
      reset_counter <= reset_counter + 8'd1;
    end else begin
      reset_counter <= reset_counter;
    end
  end
end
`endif // PALLADIUM

`ifndef WIRE_CLK
always #1 clock <= ~clock;
`endif // WIRE_CLK

SimTop sim(
  .clock(clock),
  .reset(reset),
  .difftest_logCtrl_begin(difftest_logCtrl_begin),
  .difftest_logCtrl_end(difftest_logCtrl_end),
  .difftest_logCtrl_level(difftest_logCtrl_level),
  .difftest_perfCtrl_clean(difftest_perfCtrl_clean),
  .difftest_perfCtrl_dump(difftest_perfCtrl_dump),
  .difftest_uart_out_valid(difftest_uart_out_valid),
  .difftest_uart_out_ch(difftest_uart_out_ch),
  .difftest_uart_in_valid(difftest_uart_in_valid),
  .difftest_uart_in_ch(difftest_uart_in_ch),
  .difftest_step(difftest_step)
);

assign difftest_logCtrl_level = 0;
assign difftest_perfCtrl_clean = 0;
assign difftest_perfCtrl_dump = 0;
assign difftest_uart_in_ch = 8'hff;

always @(posedge clock) begin
  if (!reset && difftest_uart_out_valid) begin
    $fwrite(32'h8000_0001, "%c", difftest_uart_out_ch);
    $fflush();
  end
end

`ifndef TB_NO_DPIC
reg [`CONFIG_DIFFTEST_STEPWIDTH - 1:0] difftest_step_delay;
always @(posedge clock) begin
  if (reset) begin
    difftest_step_delay <= 0;
  end
  else begin
    difftest_step_delay <= difftest_step;
  end
end

`ifdef CONFIG_DIFFTEST_DEFERRED_RESULT
wire simv_result;
DeferredControl deferred(
  .clock(clock),
  .reset(reset),
  .step(difftest_step_delay),
  .simv_result(simv_result)
);
`endif // CONFIG_DIFFTEST_DEFERRED_RESULT
`endif // TB_NO_DPIC

reg [63:0] n_cycles;
reg trap;
always @(posedge clock) begin
  if (reset) begin
    n_cycles <= 64'h0;
    xs_rst_en<= 1'b0;
    trap     <= 1'b0;
  end
  else if(!xs_rst_en) begin
    n_cycles <= n_cycles + 64'h1;

    // max cycles
    if (max_cycles > 0 && n_cycles >= max_cycles) begin
      $display("EXCEEDED MAX CYCLE: %d", max_cycles);
      $finish();
    end

`ifndef TB_NO_DPIC
    // difftest
    if (!n_cycles) begin
      simv_init();
      $display("simv init");
    end
`ifdef CONFIG_DIFFTEST_DEFERRED_RESULT
    else if (simv_result) begin
      $display("DIFFTEST FAILED at cycle %d", n_cycles);
      xs_rst_en <= ckpt_list_en;
    end
`else
    else if (|difftest_step_delay) begin
      // check errors
      if (trap) begin
        if (trap == 'hff && ckpt_list_en == 1'b1) begin
          $display("GCPT runing reached the maximum count point");
          xs_rst_en <= 1'b1;
        end else begin
          $display("DIFFTEST FAILED at cycle %d", n_cycles);
          $finish();
        end
      end else begin
        trap <= simv_nstep(difftest_step_delay);
      end
    end
`endif // CONFIG_DIFFTEST_DEFERRED_RESULT
`endif // TB_NO_DPIC
  end
end


always @(posedge clock)begin
  if (!reset & xs_rst_en) begin
    if (ckpt_list_en == 1'b1) begin
      if(difftest_ram_reload() == 8'd1) begin
        $display("run checkpoint end");
        $finish();
      end
    end
    else begin
      $display("not use ckpt list");
      $finish();
    end
  end
end

endmodule
