module AXI4IntrGenerator(
  input         clock,
  input         reset,
  output        auto_in_awready,
  input         auto_in_awvalid,
  input         auto_in_awid,
  input  [36:0] auto_in_awaddr,
  input  [7:0]  auto_in_awlen,
  input  [2:0]  auto_in_awsize,
  input  [1:0]  auto_in_awburst,
  input         auto_in_awlock,
  input  [3:0]  auto_in_awcache,
  input  [2:0]  auto_in_awprot,
  input  [3:0]  auto_in_awqos,
  output        auto_in_wready,
  input         auto_in_wvalid,
  input  [63:0] auto_in_wdata,
  input  [7:0]  auto_in_wstrb,
  input         auto_in_wlast,
  input         auto_in_bready,
  output        auto_in_bvalid,
  output        auto_in_bid,
  output [1:0]  auto_in_bresp,
  output        auto_in_arready,
  input         auto_in_arvalid,
  input         auto_in_arid,
  input  [36:0] auto_in_araddr,
  input  [7:0]  auto_in_arlen,
  input  [2:0]  auto_in_arsize,
  input  [1:0]  auto_in_arburst,
  input         auto_in_arlock,
  input  [3:0]  auto_in_arcache,
  input  [2:0]  auto_in_arprot,
  input  [3:0]  auto_in_arqos,
  input         auto_in_rready,
  output        auto_in_rvalid,
  output        auto_in_rid,
  output [63:0] auto_in_rdata,
  output [1:0]  auto_in_rresp,
  output        auto_in_rlast,
  output [63:0] io_extra_intrVec
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [63:0] _RAND_1015;
`endif // RANDOMIZE_REG_INIT
  wire  w_data_delay_clock; // @[Hold.scala 96:23]
  wire [31:0] w_data_delay_io_in; // @[Hold.scala 96:23]
  wire [31:0] w_data_delay_io_out; // @[Hold.scala 96:23]
  wire  delay_clock; // @[Hold.scala 96:23]
  wire [2:0] delay_io_in; // @[Hold.scala 96:23]
  wire [2:0] delay_io_out; // @[Hold.scala 96:23]
  reg [1:0] state; // @[AXI4SlaveModule.scala 95:22]
  wire  _bundleIn_0_arready_T = state == 2'h0; // @[AXI4SlaveModule.scala 153:24]
  wire  in_arready = state == 2'h0; // @[AXI4SlaveModule.scala 153:24]
  wire  in_arvalid = auto_in_arvalid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  wire  _T = in_arready & in_arvalid; // @[Decoupled.scala 50:35]
  wire  in_awready = _bundleIn_0_arready_T & ~in_arvalid; // @[AXI4SlaveModule.scala 171:35]
  wire  in_awvalid = auto_in_awvalid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  wire  _T_1 = in_awready & in_awvalid; // @[Decoupled.scala 50:35]
  wire  in_wready = state == 2'h2; // @[AXI4SlaveModule.scala 172:23]
  wire  in_wvalid = auto_in_wvalid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  wire  _T_2 = in_wready & in_wvalid; // @[Decoupled.scala 50:35]
  wire  in_bready = auto_in_bready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  wire  in_bvalid = state == 2'h3; // @[AXI4SlaveModule.scala 175:22]
  wire  _T_3 = in_bready & in_bvalid; // @[Decoupled.scala 50:35]
  wire  in_rready = auto_in_rready; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  wire  in_rvalid = state == 2'h1; // @[AXI4SlaveModule.scala 155:23]
  wire  _T_4 = in_rready & in_rvalid; // @[Decoupled.scala 50:35]
  wire [1:0] in_awburst = auto_in_awburst; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  wire [1:0] in_arburst = auto_in_arburst; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  reg [7:0] value; // @[Counter.scala 62:40]
  wire [7:0] in_arlen = auto_in_arlen; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  reg [7:0] hold_data; // @[Reg.scala 16:16]
  wire [7:0] _T_27 = _T ? in_arlen : hold_data; // @[Hold.scala 25:8]
  wire  in_rlast = value == _T_27; // @[AXI4SlaveModule.scala 133:32]
  wire  in_wlast = auto_in_wlast; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  wire [1:0] _GEN_3 = _T_2 & in_wlast ? 2'h3 : state; // @[AXI4SlaveModule.scala 112:42 113:15 95:22]
  wire [1:0] _GEN_4 = _T_3 ? 2'h0 : state; // @[AXI4SlaveModule.scala 117:24 118:15 95:22]
  wire [1:0] _GEN_5 = 2'h3 == state ? _GEN_4 : state; // @[AXI4SlaveModule.scala 97:16 95:22]
  wire [7:0] in_wstrb = auto_in_wstrb; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  reg [36:0] raddr_hold_data; // @[Reg.scala 16:16]
  wire [36:0] in_araddr = auto_in_araddr; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  wire [36:0] _GEN_10 = _T ? in_araddr : raddr_hold_data; // @[Reg.scala 16:16 17:{18,22}]
  wire [7:0] _value_T_1 = value + 8'h1; // @[Counter.scala 78:24]
  reg [36:0] waddr_hold_data; // @[Reg.scala 16:16]
  wire [36:0] in_awaddr = auto_in_awaddr; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  wire [36:0] _GEN_13 = _T_1 ? in_awaddr : waddr_hold_data; // @[Reg.scala 16:16 17:{18,22}]
  reg  bundleIn_0_bid_r; // @[Reg.scala 16:16]
  wire  in_awid = auto_in_awid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  reg  bundleIn_0_rid_r; // @[Reg.scala 16:16]
  wire  in_arid = auto_in_arid; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  reg [31:0] intrGenRegs_0; // @[AXI4IntrGenerator.scala 39:30]
  reg [31:0] intrGenRegs_1; // @[AXI4IntrGenerator.scala 39:30]
  reg [31:0] intrGenRegs_2; // @[AXI4IntrGenerator.scala 39:30]
  reg [31:0] intrGenRegs_3; // @[AXI4IntrGenerator.scala 39:30]
  reg [31:0] intrGenRegs_4; // @[AXI4IntrGenerator.scala 39:30]
  reg [31:0] intrGenRegs_5; // @[AXI4IntrGenerator.scala 39:30]
  reg [31:0] intrGenRegs_6; // @[AXI4IntrGenerator.scala 39:30]
  reg [63:0] randomPosition_lfsr; // @[LFSR64.scala 25:23]
  wire  randomPosition_xor = randomPosition_lfsr[0] ^ randomPosition_lfsr[1] ^ randomPosition_lfsr[3] ^
    randomPosition_lfsr[4]; // @[LFSR64.scala 26:43]
  wire [63:0] _randomPosition_lfsr_T_2 = {randomPosition_xor,randomPosition_lfsr[63:1]}; // @[Cat.scala 31:58]
  wire [5:0] randomPosition = randomPosition_lfsr[5:0]; // @[AXI4IntrGenerator.scala 50:34]
  wire [31:0] _GEN_20 = randomPosition[5] ? intrGenRegs_3 : intrGenRegs_2; // @[AXI4IntrGenerator.scala 51:{85,85}]
  wire [31:0] _randomCondition_T_3 = _GEN_20 >> randomPosition[4:0]; // @[AXI4IntrGenerator.scala 51:85]
  wire  randomCondition = intrGenRegs_5 == intrGenRegs_6 & _randomCondition_T_3[0]; // @[AXI4IntrGenerator.scala 51:53]
  wire [31:0] _intrGenRegs_5_T_1 = intrGenRegs_5 + 32'h1; // @[AXI4IntrGenerator.scala 52:32]
  wire [31:0] _intrGenRegs_T_2 = 32'h1 << randomPosition[4:0]; // @[OneHot.scala 57:35]
  wire [31:0] _GEN_22 = randomPosition[5] ? intrGenRegs_1 : intrGenRegs_0; // @[AXI4IntrGenerator.scala 54:{68,68}]
  wire [31:0] _intrGenRegs_T_3 = _GEN_22 | _intrGenRegs_T_2; // @[AXI4IntrGenerator.scala 54:68]
  wire [31:0] _GEN_23 = ~randomPosition[5] ? _intrGenRegs_T_3 : intrGenRegs_0; // @[AXI4IntrGenerator.scala 39:30 54:{38,38}]
  wire [31:0] _GEN_24 = randomPosition[5] ? _intrGenRegs_T_3 : intrGenRegs_1; // @[AXI4IntrGenerator.scala 39:30 54:{38,38}]
  wire [1:0] _GEN_76 = {{1'd0}, randomPosition[5]}; // @[AXI4IntrGenerator.scala 39:30 54:{38,38}]
  wire [31:0] _GEN_25 = 2'h2 == _GEN_76 ? _intrGenRegs_T_3 : intrGenRegs_2; // @[AXI4IntrGenerator.scala 39:30 54:{38,38}]
  wire [31:0] _GEN_26 = 2'h3 == _GEN_76 ? _intrGenRegs_T_3 : intrGenRegs_3; // @[AXI4IntrGenerator.scala 39:30 54:{38,38}]
  wire [2:0] _GEN_78 = {{2'd0}, randomPosition[5]}; // @[AXI4IntrGenerator.scala 39:30 54:{38,38}]
  wire [31:0] _GEN_27 = 3'h4 == _GEN_78 ? _intrGenRegs_T_3 : intrGenRegs_4; // @[AXI4IntrGenerator.scala 39:30 54:{38,38}]
  wire [31:0] _GEN_28 = 3'h5 == _GEN_78 ? _intrGenRegs_T_3 : _intrGenRegs_5_T_1; // @[AXI4IntrGenerator.scala 52:17 54:{38,38}]
  wire [31:0] _GEN_29 = 3'h6 == _GEN_78 ? _intrGenRegs_T_3 : intrGenRegs_6; // @[AXI4IntrGenerator.scala 39:30 54:{38,38}]
  wire [31:0] _GEN_31 = randomCondition ? _GEN_23 : intrGenRegs_0; // @[AXI4IntrGenerator.scala 53:28 39:30]
  wire [31:0] _GEN_32 = randomCondition ? _GEN_24 : intrGenRegs_1; // @[AXI4IntrGenerator.scala 53:28 39:30]
  wire [31:0] _GEN_33 = randomCondition ? _GEN_25 : intrGenRegs_2; // @[AXI4IntrGenerator.scala 53:28 39:30]
  wire [31:0] _GEN_34 = randomCondition ? _GEN_26 : intrGenRegs_3; // @[AXI4IntrGenerator.scala 53:28 39:30]
  wire [31:0] _GEN_35 = randomCondition ? _GEN_27 : intrGenRegs_4; // @[AXI4IntrGenerator.scala 53:28 39:30]
  wire [31:0] _GEN_36 = randomCondition ? _GEN_28 : _intrGenRegs_5_T_1; // @[AXI4IntrGenerator.scala 52:17 53:28]
  wire [31:0] _GEN_37 = randomCondition ? _GEN_29 : intrGenRegs_6; // @[AXI4IntrGenerator.scala 53:28 39:30]
  wire [63:0] in_wdata = auto_in_wdata; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  wire  w_fire = _T_2 & in_wdata != 64'h0; // @[AXI4IntrGenerator.scala 61:28]
  reg  REG; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_1; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_2; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_3; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_4; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_5; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_6; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_7; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_8; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_9; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_10; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_11; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_12; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_13; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_14; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_15; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_16; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_17; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_18; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_19; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_20; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_21; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_22; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_23; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_24; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_25; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_26; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_27; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_28; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_29; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_30; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_31; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_32; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_33; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_34; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_35; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_36; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_37; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_38; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_39; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_40; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_41; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_42; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_43; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_44; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_45; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_46; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_47; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_48; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_49; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_50; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_51; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_52; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_53; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_54; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_55; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_56; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_57; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_58; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_59; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_60; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_61; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_62; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_63; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_64; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_65; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_66; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_67; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_68; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_69; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_70; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_71; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_72; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_73; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_74; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_75; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_76; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_77; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_78; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_79; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_80; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_81; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_82; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_83; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_84; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_85; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_86; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_87; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_88; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_89; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_90; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_91; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_92; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_93; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_94; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_95; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_96; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_97; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_98; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_99; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_100; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_101; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_102; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_103; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_104; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_105; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_106; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_107; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_108; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_109; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_110; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_111; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_112; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_113; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_114; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_115; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_116; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_117; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_118; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_119; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_120; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_121; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_122; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_123; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_124; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_125; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_126; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_127; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_128; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_129; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_130; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_131; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_132; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_133; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_134; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_135; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_136; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_137; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_138; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_139; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_140; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_141; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_142; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_143; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_144; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_145; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_146; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_147; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_148; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_149; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_150; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_151; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_152; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_153; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_154; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_155; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_156; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_157; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_158; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_159; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_160; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_161; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_162; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_163; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_164; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_165; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_166; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_167; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_168; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_169; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_170; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_171; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_172; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_173; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_174; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_175; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_176; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_177; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_178; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_179; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_180; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_181; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_182; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_183; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_184; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_185; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_186; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_187; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_188; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_189; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_190; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_191; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_192; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_193; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_194; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_195; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_196; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_197; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_198; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_199; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_200; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_201; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_202; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_203; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_204; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_205; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_206; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_207; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_208; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_209; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_210; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_211; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_212; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_213; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_214; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_215; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_216; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_217; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_218; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_219; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_220; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_221; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_222; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_223; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_224; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_225; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_226; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_227; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_228; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_229; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_230; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_231; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_232; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_233; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_234; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_235; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_236; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_237; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_238; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_239; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_240; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_241; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_242; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_243; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_244; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_245; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_246; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_247; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_248; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_249; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_250; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_251; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_252; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_253; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_254; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_255; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_256; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_257; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_258; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_259; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_260; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_261; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_262; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_263; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_264; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_265; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_266; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_267; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_268; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_269; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_270; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_271; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_272; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_273; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_274; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_275; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_276; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_277; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_278; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_279; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_280; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_281; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_282; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_283; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_284; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_285; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_286; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_287; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_288; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_289; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_290; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_291; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_292; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_293; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_294; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_295; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_296; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_297; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_298; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_299; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_300; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_301; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_302; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_303; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_304; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_305; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_306; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_307; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_308; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_309; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_310; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_311; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_312; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_313; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_314; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_315; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_316; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_317; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_318; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_319; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_320; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_321; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_322; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_323; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_324; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_325; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_326; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_327; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_328; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_329; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_330; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_331; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_332; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_333; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_334; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_335; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_336; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_337; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_338; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_339; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_340; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_341; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_342; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_343; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_344; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_345; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_346; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_347; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_348; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_349; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_350; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_351; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_352; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_353; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_354; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_355; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_356; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_357; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_358; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_359; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_360; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_361; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_362; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_363; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_364; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_365; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_366; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_367; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_368; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_369; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_370; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_371; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_372; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_373; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_374; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_375; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_376; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_377; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_378; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_379; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_380; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_381; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_382; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_383; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_384; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_385; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_386; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_387; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_388; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_389; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_390; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_391; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_392; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_393; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_394; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_395; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_396; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_397; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_398; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_399; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_400; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_401; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_402; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_403; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_404; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_405; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_406; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_407; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_408; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_409; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_410; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_411; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_412; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_413; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_414; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_415; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_416; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_417; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_418; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_419; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_420; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_421; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_422; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_423; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_424; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_425; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_426; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_427; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_428; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_429; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_430; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_431; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_432; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_433; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_434; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_435; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_436; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_437; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_438; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_439; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_440; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_441; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_442; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_443; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_444; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_445; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_446; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_447; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_448; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_449; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_450; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_451; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_452; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_453; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_454; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_455; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_456; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_457; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_458; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_459; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_460; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_461; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_462; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_463; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_464; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_465; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_466; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_467; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_468; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_469; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_470; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_471; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_472; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_473; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_474; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_475; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_476; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_477; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_478; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_479; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_480; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_481; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_482; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_483; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_484; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_485; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_486; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_487; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_488; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_489; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_490; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_491; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_492; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_493; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_494; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_495; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_496; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_497; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_498; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_499; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_500; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_501; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_502; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_503; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_504; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_505; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_506; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_507; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_508; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_509; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_510; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_511; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_512; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_513; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_514; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_515; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_516; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_517; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_518; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_519; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_520; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_521; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_522; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_523; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_524; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_525; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_526; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_527; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_528; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_529; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_530; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_531; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_532; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_533; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_534; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_535; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_536; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_537; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_538; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_539; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_540; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_541; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_542; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_543; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_544; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_545; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_546; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_547; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_548; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_549; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_550; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_551; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_552; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_553; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_554; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_555; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_556; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_557; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_558; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_559; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_560; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_561; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_562; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_563; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_564; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_565; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_566; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_567; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_568; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_569; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_570; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_571; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_572; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_573; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_574; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_575; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_576; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_577; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_578; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_579; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_580; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_581; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_582; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_583; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_584; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_585; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_586; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_587; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_588; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_589; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_590; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_591; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_592; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_593; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_594; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_595; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_596; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_597; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_598; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_599; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_600; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_601; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_602; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_603; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_604; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_605; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_606; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_607; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_608; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_609; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_610; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_611; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_612; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_613; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_614; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_615; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_616; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_617; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_618; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_619; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_620; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_621; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_622; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_623; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_624; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_625; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_626; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_627; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_628; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_629; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_630; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_631; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_632; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_633; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_634; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_635; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_636; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_637; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_638; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_639; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_640; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_641; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_642; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_643; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_644; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_645; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_646; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_647; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_648; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_649; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_650; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_651; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_652; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_653; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_654; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_655; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_656; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_657; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_658; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_659; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_660; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_661; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_662; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_663; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_664; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_665; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_666; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_667; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_668; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_669; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_670; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_671; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_672; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_673; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_674; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_675; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_676; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_677; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_678; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_679; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_680; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_681; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_682; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_683; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_684; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_685; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_686; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_687; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_688; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_689; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_690; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_691; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_692; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_693; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_694; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_695; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_696; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_697; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_698; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_699; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_700; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_701; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_702; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_703; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_704; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_705; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_706; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_707; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_708; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_709; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_710; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_711; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_712; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_713; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_714; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_715; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_716; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_717; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_718; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_719; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_720; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_721; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_722; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_723; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_724; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_725; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_726; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_727; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_728; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_729; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_730; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_731; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_732; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_733; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_734; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_735; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_736; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_737; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_738; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_739; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_740; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_741; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_742; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_743; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_744; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_745; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_746; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_747; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_748; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_749; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_750; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_751; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_752; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_753; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_754; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_755; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_756; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_757; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_758; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_759; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_760; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_761; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_762; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_763; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_764; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_765; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_766; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_767; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_768; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_769; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_770; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_771; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_772; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_773; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_774; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_775; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_776; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_777; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_778; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_779; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_780; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_781; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_782; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_783; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_784; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_785; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_786; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_787; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_788; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_789; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_790; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_791; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_792; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_793; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_794; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_795; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_796; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_797; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_798; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_799; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_800; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_801; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_802; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_803; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_804; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_805; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_806; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_807; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_808; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_809; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_810; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_811; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_812; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_813; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_814; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_815; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_816; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_817; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_818; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_819; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_820; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_821; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_822; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_823; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_824; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_825; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_826; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_827; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_828; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_829; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_830; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_831; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_832; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_833; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_834; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_835; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_836; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_837; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_838; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_839; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_840; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_841; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_842; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_843; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_844; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_845; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_846; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_847; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_848; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_849; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_850; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_851; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_852; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_853; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_854; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_855; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_856; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_857; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_858; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_859; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_860; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_861; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_862; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_863; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_864; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_865; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_866; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_867; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_868; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_869; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_870; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_871; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_872; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_873; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_874; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_875; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_876; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_877; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_878; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_879; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_880; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_881; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_882; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_883; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_884; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_885; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_886; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_887; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_888; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_889; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_890; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_891; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_892; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_893; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_894; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_895; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_896; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_897; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_898; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_899; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_900; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_901; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_902; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_903; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_904; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_905; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_906; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_907; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_908; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_909; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_910; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_911; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_912; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_913; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_914; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_915; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_916; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_917; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_918; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_919; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_920; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_921; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_922; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_923; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_924; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_925; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_926; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_927; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_928; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_929; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_930; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_931; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_932; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_933; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_934; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_935; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_936; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_937; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_938; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_939; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_940; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_941; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_942; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_943; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_944; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_945; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_946; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_947; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_948; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_949; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_950; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_951; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_952; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_953; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_954; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_955; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_956; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_957; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_958; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_959; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_960; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_961; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_962; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_963; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_964; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_965; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_966; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_967; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_968; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_969; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_970; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_971; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_972; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_973; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_974; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_975; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_976; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_977; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_978; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_979; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_980; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_981; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_982; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_983; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_984; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_985; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_986; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_987; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_988; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_989; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_990; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_991; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_992; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_993; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_994; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_995; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_996; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_997; // @[AXI4IntrGenerator.scala 63:23]
  reg  REG_998; // @[AXI4IntrGenerator.scala 63:23]
  reg  w_fire_1; // @[AXI4IntrGenerator.scala 63:23]
  wire [31:0] _intrGenRegs_delay_io_out = w_data_delay_io_out; // @[AXI4IntrGenerator.scala 67:{53,53}]
  wire [31:0] _GEN_39 = 3'h0 == delay_io_out ? _intrGenRegs_delay_io_out : _GEN_31; // @[AXI4IntrGenerator.scala 67:{53,53}]
  wire [31:0] _GEN_40 = 3'h1 == delay_io_out ? _intrGenRegs_delay_io_out : _GEN_32; // @[AXI4IntrGenerator.scala 67:{53,53}]
  wire [31:0] _GEN_41 = 3'h2 == delay_io_out ? _intrGenRegs_delay_io_out : _GEN_33; // @[AXI4IntrGenerator.scala 67:{53,53}]
  wire [31:0] _GEN_42 = 3'h3 == delay_io_out ? _intrGenRegs_delay_io_out : _GEN_34; // @[AXI4IntrGenerator.scala 67:{53,53}]
  wire [31:0] _GEN_43 = 3'h4 == delay_io_out ? _intrGenRegs_delay_io_out : _GEN_35; // @[AXI4IntrGenerator.scala 67:{53,53}]
  wire [31:0] _GEN_44 = 3'h5 == delay_io_out ? _intrGenRegs_delay_io_out : _GEN_36; // @[AXI4IntrGenerator.scala 67:{53,53}]
  wire [31:0] _GEN_45 = 3'h6 == delay_io_out ? _intrGenRegs_delay_io_out : _GEN_37; // @[AXI4IntrGenerator.scala 67:{53,53}]
  wire [31:0] _GEN_47 = w_fire_1 ? _GEN_39 : _GEN_31; // @[AXI4IntrGenerator.scala 66:19]
  wire [31:0] _GEN_48 = w_fire_1 ? _GEN_40 : _GEN_32; // @[AXI4IntrGenerator.scala 66:19]
  wire [31:0] _GEN_49 = w_fire_1 ? _GEN_41 : _GEN_33; // @[AXI4IntrGenerator.scala 66:19]
  wire [31:0] _GEN_50 = w_fire_1 ? _GEN_42 : _GEN_34; // @[AXI4IntrGenerator.scala 66:19]
  wire [31:0] _GEN_51 = w_fire_1 ? _GEN_43 : _GEN_35; // @[AXI4IntrGenerator.scala 66:19]
  wire [31:0] _GEN_52 = w_fire_1 ? _GEN_44 : _GEN_36; // @[AXI4IntrGenerator.scala 66:19]
  wire [31:0] _GEN_53 = w_fire_1 ? _GEN_45 : _GEN_37; // @[AXI4IntrGenerator.scala 66:19]
  wire  _T_47 = _T_2 & in_wdata == 64'h0; // @[AXI4IntrGenerator.scala 70:21]
  wire [31:0] _GEN_61 = 3'h6 == _GEN_13[4:2] ? 32'h0 : _GEN_53; // @[AXI4IntrGenerator.scala 71:{32,32}]
  wire [31:0] _GEN_69 = _T_2 & in_wdata == 64'h0 ? _GEN_61 : _GEN_53; // @[AXI4IntrGenerator.scala 70:48]
  reg [63:0] intrGenRegs_6_lfsr; // @[LFSR64.scala 25:23]
  wire  intrGenRegs_6_xor = intrGenRegs_6_lfsr[0] ^ intrGenRegs_6_lfsr[1] ^ intrGenRegs_6_lfsr[3] ^ intrGenRegs_6_lfsr[4
    ]; // @[LFSR64.scala 26:43]
  wire [63:0] _intrGenRegs_6_lfsr_T_2 = {intrGenRegs_6_xor,intrGenRegs_6_lfsr[63:1]}; // @[Cat.scala 31:58]
  wire [63:0] _GEN_82 = {{32'd0}, intrGenRegs_4}; // @[AXI4IntrGenerator.scala 75:29]
  wire [63:0] _intrGenRegs_6_T = intrGenRegs_6_lfsr & _GEN_82; // @[AXI4IntrGenerator.scala 75:29]
  wire [63:0] _GEN_72 = _T_47 | w_fire_1 ? _intrGenRegs_6_T : {{32'd0}, _GEN_69}; // @[AXI4IntrGenerator.scala 74:58 75:17]
  wire [31:0] _GEN_75 = _GEN_10[0] ? intrGenRegs_1 : intrGenRegs_0; // @[AXI4IntrGenerator.scala 79:{20,20}]
  wire [7:0] in_awlen = auto_in_awlen; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  wire [2:0] in_awsize = auto_in_awsize; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  wire  in_awlock = auto_in_awlock; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  wire [3:0] in_awcache = auto_in_awcache; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  wire [2:0] in_awprot = auto_in_awprot; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  wire [3:0] in_awqos = auto_in_awqos; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  wire  in_bid = bundleIn_0_bid_r; // @[Nodes.scala 1210:84 AXI4SlaveModule.scala 177:16]
  wire [1:0] in_bresp = 2'h0; // @[Nodes.scala 1210:84 AXI4SlaveModule.scala 174:18]
  wire [2:0] in_arsize = auto_in_arsize; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  wire  in_arlock = auto_in_arlock; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  wire [3:0] in_arcache = auto_in_arcache; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  wire [2:0] in_arprot = auto_in_arprot; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  wire [3:0] in_arqos = auto_in_arqos; // @[Nodes.scala 1210:84 LazyModule.scala 309:16]
  wire  in_rid = bundleIn_0_rid_r; // @[Nodes.scala 1210:84 AXI4SlaveModule.scala 179:16]
  wire [63:0] in_rdata = {{32'd0}, _GEN_75}; // @[Nodes.scala 1210:84 AXI4IntrGenerator.scala 79:20]
  wire [1:0] in_rresp = 2'h0; // @[Nodes.scala 1210:84 AXI4SlaveModule.scala 154:18]
  wire [63:0] _GEN_83 = reset ? 64'h0 : _GEN_72; // @[AXI4IntrGenerator.scala 39:{30,30}]
  DelayN_36 w_data_delay ( // @[Hold.scala 96:23]
    .clock(w_data_delay_clock),
    .io_in(w_data_delay_io_in),
    .io_out(w_data_delay_io_out)
  );
  DelayN_37 delay ( // @[Hold.scala 96:23]
    .clock(delay_clock),
    .io_in(delay_io_in),
    .io_out(delay_io_out)
  );
  assign auto_in_awready = in_awready; // @[LazyModule.scala 309:16]
  assign auto_in_wready = in_wready; // @[LazyModule.scala 309:16]
  assign auto_in_bvalid = in_bvalid; // @[LazyModule.scala 309:16]
  assign auto_in_bid = in_bid; // @[LazyModule.scala 309:16]
  assign auto_in_bresp = in_bresp; // @[LazyModule.scala 309:16]
  assign auto_in_arready = in_arready; // @[LazyModule.scala 309:16]
  assign auto_in_rvalid = in_rvalid; // @[LazyModule.scala 309:16]
  assign auto_in_rid = in_rid; // @[LazyModule.scala 309:16]
  assign auto_in_rdata = in_rdata; // @[LazyModule.scala 309:16]
  assign auto_in_rresp = in_bresp; // @[LazyModule.scala 309:16]
  assign auto_in_rlast = in_rlast; // @[LazyModule.scala 309:16]
  assign io_extra_intrVec = {intrGenRegs_1,intrGenRegs_0}; // @[Cat.scala 31:58]
  assign w_data_delay_clock = clock;
  assign w_data_delay_io_in = in_wdata[31:0]; // @[AXI4IntrGenerator.scala 65:39]
  assign delay_clock = clock;
  assign delay_io_in = _GEN_13[4:2]; // @[AXI4IntrGenerator.scala 67:31]
  always @(posedge clock) begin
    if (reset) begin // @[AXI4SlaveModule.scala 95:22]
      state <= 2'h0; // @[AXI4SlaveModule.scala 95:22]
    end else if (2'h0 == state) begin // @[AXI4SlaveModule.scala 97:16]
      if (_T_1) begin // @[AXI4SlaveModule.scala 102:25]
        state <= 2'h2; // @[AXI4SlaveModule.scala 103:15]
      end else if (_T) begin // @[AXI4SlaveModule.scala 99:25]
        state <= 2'h1; // @[AXI4SlaveModule.scala 100:15]
      end
    end else if (2'h1 == state) begin // @[AXI4SlaveModule.scala 97:16]
      if (_T_4 & in_rlast) begin // @[AXI4SlaveModule.scala 107:42]
        state <= 2'h0; // @[AXI4SlaveModule.scala 108:15]
      end
    end else if (2'h2 == state) begin // @[AXI4SlaveModule.scala 97:16]
      state <= _GEN_3;
    end else begin
      state <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      value <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_4) begin // @[AXI4SlaveModule.scala 135:23]
      if (in_rlast) begin // @[AXI4SlaveModule.scala 137:28]
        value <= 8'h0; // @[AXI4SlaveModule.scala 138:17]
      end else begin
        value <= _value_T_1; // @[Counter.scala 78:15]
      end
    end
    if (_T) begin // @[Reg.scala 17:18]
      hold_data <= in_arlen; // @[Reg.scala 17:22]
    end
    if (_T) begin // @[Reg.scala 17:18]
      raddr_hold_data <= in_araddr; // @[Reg.scala 17:22]
    end
    if (_T_1) begin // @[Reg.scala 17:18]
      waddr_hold_data <= in_awaddr; // @[Reg.scala 17:22]
    end
    if (_T_1) begin // @[Reg.scala 17:18]
      bundleIn_0_bid_r <= in_awid; // @[Reg.scala 17:22]
    end
    if (_T) begin // @[Reg.scala 17:18]
      bundleIn_0_rid_r <= in_arid; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 39:30]
      intrGenRegs_0 <= 32'h0; // @[AXI4IntrGenerator.scala 39:30]
    end else if (_T_2 & in_wdata == 64'h0) begin // @[AXI4IntrGenerator.scala 70:48]
      if (3'h0 == _GEN_13[4:2]) begin // @[AXI4IntrGenerator.scala 71:32]
        intrGenRegs_0 <= 32'h0; // @[AXI4IntrGenerator.scala 71:32]
      end else begin
        intrGenRegs_0 <= _GEN_47;
      end
    end else begin
      intrGenRegs_0 <= _GEN_47;
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 39:30]
      intrGenRegs_1 <= 32'h0; // @[AXI4IntrGenerator.scala 39:30]
    end else if (_T_2 & in_wdata == 64'h0) begin // @[AXI4IntrGenerator.scala 70:48]
      if (3'h1 == _GEN_13[4:2]) begin // @[AXI4IntrGenerator.scala 71:32]
        intrGenRegs_1 <= 32'h0; // @[AXI4IntrGenerator.scala 71:32]
      end else begin
        intrGenRegs_1 <= _GEN_48;
      end
    end else begin
      intrGenRegs_1 <= _GEN_48;
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 39:30]
      intrGenRegs_2 <= 32'h0; // @[AXI4IntrGenerator.scala 39:30]
    end else if (_T_2 & in_wdata == 64'h0) begin // @[AXI4IntrGenerator.scala 70:48]
      if (3'h2 == _GEN_13[4:2]) begin // @[AXI4IntrGenerator.scala 71:32]
        intrGenRegs_2 <= 32'h0; // @[AXI4IntrGenerator.scala 71:32]
      end else begin
        intrGenRegs_2 <= _GEN_49;
      end
    end else begin
      intrGenRegs_2 <= _GEN_49;
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 39:30]
      intrGenRegs_3 <= 32'h0; // @[AXI4IntrGenerator.scala 39:30]
    end else if (_T_2 & in_wdata == 64'h0) begin // @[AXI4IntrGenerator.scala 70:48]
      if (3'h3 == _GEN_13[4:2]) begin // @[AXI4IntrGenerator.scala 71:32]
        intrGenRegs_3 <= 32'h0; // @[AXI4IntrGenerator.scala 71:32]
      end else begin
        intrGenRegs_3 <= _GEN_50;
      end
    end else begin
      intrGenRegs_3 <= _GEN_50;
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 39:30]
      intrGenRegs_4 <= 32'h0; // @[AXI4IntrGenerator.scala 39:30]
    end else if (_T_2 & in_wdata == 64'h0) begin // @[AXI4IntrGenerator.scala 70:48]
      if (3'h4 == _GEN_13[4:2]) begin // @[AXI4IntrGenerator.scala 71:32]
        intrGenRegs_4 <= 32'h0; // @[AXI4IntrGenerator.scala 71:32]
      end else begin
        intrGenRegs_4 <= _GEN_51;
      end
    end else begin
      intrGenRegs_4 <= _GEN_51;
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 39:30]
      intrGenRegs_5 <= 32'h0; // @[AXI4IntrGenerator.scala 39:30]
    end else if (_T_47 | w_fire_1) begin // @[AXI4IntrGenerator.scala 74:58]
      intrGenRegs_5 <= 32'h0; // @[AXI4IntrGenerator.scala 76:19]
    end else if (_T_2 & in_wdata == 64'h0) begin // @[AXI4IntrGenerator.scala 70:48]
      if (3'h5 == _GEN_13[4:2]) begin // @[AXI4IntrGenerator.scala 71:32]
        intrGenRegs_5 <= 32'h0; // @[AXI4IntrGenerator.scala 71:32]
      end else begin
        intrGenRegs_5 <= _GEN_52;
      end
    end else begin
      intrGenRegs_5 <= _GEN_52;
    end
    intrGenRegs_6 <= _GEN_83[31:0]; // @[AXI4IntrGenerator.scala 39:{30,30}]
    if (reset) begin // @[LFSR64.scala 25:23]
      randomPosition_lfsr <= 64'h1234567887654321; // @[LFSR64.scala 25:23]
    end else if (randomPosition_lfsr == 64'h0) begin // @[LFSR64.scala 28:18]
      randomPosition_lfsr <= 64'h1;
    end else begin
      randomPosition_lfsr <= _randomPosition_lfsr_T_2;
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG <= w_fire; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_1 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_1 <= REG; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_2 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_2 <= REG_1; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_3 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_3 <= REG_2; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_4 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_4 <= REG_3; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_5 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_5 <= REG_4; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_6 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_6 <= REG_5; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_7 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_7 <= REG_6; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_8 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_8 <= REG_7; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_9 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_9 <= REG_8; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_10 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_10 <= REG_9; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_11 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_11 <= REG_10; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_12 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_12 <= REG_11; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_13 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_13 <= REG_12; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_14 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_14 <= REG_13; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_15 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_15 <= REG_14; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_16 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_16 <= REG_15; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_17 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_17 <= REG_16; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_18 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_18 <= REG_17; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_19 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_19 <= REG_18; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_20 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_20 <= REG_19; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_21 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_21 <= REG_20; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_22 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_22 <= REG_21; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_23 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_23 <= REG_22; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_24 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_24 <= REG_23; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_25 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_25 <= REG_24; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_26 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_26 <= REG_25; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_27 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_27 <= REG_26; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_28 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_28 <= REG_27; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_29 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_29 <= REG_28; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_30 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_30 <= REG_29; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_31 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_31 <= REG_30; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_32 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_32 <= REG_31; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_33 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_33 <= REG_32; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_34 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_34 <= REG_33; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_35 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_35 <= REG_34; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_36 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_36 <= REG_35; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_37 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_37 <= REG_36; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_38 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_38 <= REG_37; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_39 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_39 <= REG_38; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_40 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_40 <= REG_39; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_41 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_41 <= REG_40; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_42 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_42 <= REG_41; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_43 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_43 <= REG_42; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_44 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_44 <= REG_43; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_45 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_45 <= REG_44; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_46 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_46 <= REG_45; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_47 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_47 <= REG_46; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_48 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_48 <= REG_47; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_49 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_49 <= REG_48; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_50 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_50 <= REG_49; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_51 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_51 <= REG_50; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_52 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_52 <= REG_51; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_53 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_53 <= REG_52; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_54 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_54 <= REG_53; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_55 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_55 <= REG_54; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_56 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_56 <= REG_55; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_57 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_57 <= REG_56; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_58 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_58 <= REG_57; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_59 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_59 <= REG_58; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_60 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_60 <= REG_59; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_61 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_61 <= REG_60; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_62 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_62 <= REG_61; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_63 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_63 <= REG_62; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_64 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_64 <= REG_63; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_65 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_65 <= REG_64; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_66 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_66 <= REG_65; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_67 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_67 <= REG_66; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_68 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_68 <= REG_67; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_69 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_69 <= REG_68; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_70 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_70 <= REG_69; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_71 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_71 <= REG_70; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_72 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_72 <= REG_71; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_73 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_73 <= REG_72; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_74 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_74 <= REG_73; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_75 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_75 <= REG_74; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_76 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_76 <= REG_75; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_77 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_77 <= REG_76; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_78 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_78 <= REG_77; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_79 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_79 <= REG_78; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_80 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_80 <= REG_79; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_81 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_81 <= REG_80; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_82 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_82 <= REG_81; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_83 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_83 <= REG_82; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_84 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_84 <= REG_83; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_85 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_85 <= REG_84; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_86 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_86 <= REG_85; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_87 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_87 <= REG_86; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_88 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_88 <= REG_87; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_89 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_89 <= REG_88; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_90 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_90 <= REG_89; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_91 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_91 <= REG_90; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_92 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_92 <= REG_91; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_93 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_93 <= REG_92; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_94 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_94 <= REG_93; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_95 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_95 <= REG_94; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_96 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_96 <= REG_95; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_97 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_97 <= REG_96; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_98 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_98 <= REG_97; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_99 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_99 <= REG_98; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_100 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_100 <= REG_99; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_101 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_101 <= REG_100; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_102 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_102 <= REG_101; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_103 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_103 <= REG_102; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_104 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_104 <= REG_103; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_105 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_105 <= REG_104; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_106 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_106 <= REG_105; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_107 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_107 <= REG_106; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_108 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_108 <= REG_107; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_109 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_109 <= REG_108; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_110 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_110 <= REG_109; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_111 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_111 <= REG_110; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_112 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_112 <= REG_111; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_113 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_113 <= REG_112; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_114 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_114 <= REG_113; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_115 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_115 <= REG_114; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_116 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_116 <= REG_115; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_117 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_117 <= REG_116; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_118 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_118 <= REG_117; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_119 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_119 <= REG_118; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_120 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_120 <= REG_119; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_121 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_121 <= REG_120; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_122 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_122 <= REG_121; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_123 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_123 <= REG_122; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_124 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_124 <= REG_123; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_125 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_125 <= REG_124; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_126 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_126 <= REG_125; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_127 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_127 <= REG_126; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_128 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_128 <= REG_127; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_129 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_129 <= REG_128; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_130 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_130 <= REG_129; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_131 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_131 <= REG_130; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_132 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_132 <= REG_131; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_133 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_133 <= REG_132; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_134 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_134 <= REG_133; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_135 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_135 <= REG_134; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_136 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_136 <= REG_135; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_137 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_137 <= REG_136; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_138 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_138 <= REG_137; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_139 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_139 <= REG_138; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_140 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_140 <= REG_139; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_141 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_141 <= REG_140; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_142 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_142 <= REG_141; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_143 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_143 <= REG_142; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_144 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_144 <= REG_143; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_145 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_145 <= REG_144; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_146 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_146 <= REG_145; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_147 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_147 <= REG_146; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_148 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_148 <= REG_147; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_149 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_149 <= REG_148; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_150 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_150 <= REG_149; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_151 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_151 <= REG_150; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_152 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_152 <= REG_151; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_153 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_153 <= REG_152; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_154 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_154 <= REG_153; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_155 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_155 <= REG_154; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_156 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_156 <= REG_155; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_157 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_157 <= REG_156; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_158 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_158 <= REG_157; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_159 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_159 <= REG_158; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_160 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_160 <= REG_159; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_161 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_161 <= REG_160; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_162 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_162 <= REG_161; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_163 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_163 <= REG_162; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_164 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_164 <= REG_163; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_165 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_165 <= REG_164; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_166 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_166 <= REG_165; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_167 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_167 <= REG_166; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_168 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_168 <= REG_167; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_169 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_169 <= REG_168; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_170 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_170 <= REG_169; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_171 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_171 <= REG_170; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_172 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_172 <= REG_171; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_173 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_173 <= REG_172; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_174 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_174 <= REG_173; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_175 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_175 <= REG_174; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_176 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_176 <= REG_175; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_177 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_177 <= REG_176; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_178 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_178 <= REG_177; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_179 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_179 <= REG_178; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_180 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_180 <= REG_179; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_181 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_181 <= REG_180; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_182 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_182 <= REG_181; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_183 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_183 <= REG_182; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_184 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_184 <= REG_183; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_185 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_185 <= REG_184; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_186 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_186 <= REG_185; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_187 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_187 <= REG_186; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_188 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_188 <= REG_187; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_189 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_189 <= REG_188; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_190 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_190 <= REG_189; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_191 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_191 <= REG_190; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_192 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_192 <= REG_191; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_193 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_193 <= REG_192; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_194 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_194 <= REG_193; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_195 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_195 <= REG_194; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_196 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_196 <= REG_195; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_197 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_197 <= REG_196; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_198 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_198 <= REG_197; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_199 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_199 <= REG_198; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_200 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_200 <= REG_199; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_201 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_201 <= REG_200; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_202 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_202 <= REG_201; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_203 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_203 <= REG_202; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_204 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_204 <= REG_203; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_205 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_205 <= REG_204; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_206 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_206 <= REG_205; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_207 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_207 <= REG_206; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_208 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_208 <= REG_207; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_209 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_209 <= REG_208; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_210 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_210 <= REG_209; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_211 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_211 <= REG_210; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_212 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_212 <= REG_211; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_213 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_213 <= REG_212; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_214 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_214 <= REG_213; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_215 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_215 <= REG_214; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_216 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_216 <= REG_215; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_217 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_217 <= REG_216; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_218 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_218 <= REG_217; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_219 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_219 <= REG_218; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_220 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_220 <= REG_219; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_221 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_221 <= REG_220; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_222 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_222 <= REG_221; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_223 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_223 <= REG_222; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_224 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_224 <= REG_223; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_225 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_225 <= REG_224; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_226 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_226 <= REG_225; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_227 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_227 <= REG_226; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_228 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_228 <= REG_227; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_229 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_229 <= REG_228; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_230 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_230 <= REG_229; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_231 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_231 <= REG_230; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_232 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_232 <= REG_231; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_233 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_233 <= REG_232; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_234 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_234 <= REG_233; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_235 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_235 <= REG_234; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_236 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_236 <= REG_235; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_237 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_237 <= REG_236; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_238 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_238 <= REG_237; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_239 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_239 <= REG_238; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_240 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_240 <= REG_239; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_241 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_241 <= REG_240; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_242 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_242 <= REG_241; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_243 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_243 <= REG_242; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_244 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_244 <= REG_243; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_245 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_245 <= REG_244; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_246 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_246 <= REG_245; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_247 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_247 <= REG_246; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_248 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_248 <= REG_247; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_249 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_249 <= REG_248; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_250 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_250 <= REG_249; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_251 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_251 <= REG_250; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_252 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_252 <= REG_251; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_253 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_253 <= REG_252; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_254 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_254 <= REG_253; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_255 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_255 <= REG_254; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_256 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_256 <= REG_255; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_257 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_257 <= REG_256; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_258 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_258 <= REG_257; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_259 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_259 <= REG_258; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_260 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_260 <= REG_259; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_261 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_261 <= REG_260; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_262 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_262 <= REG_261; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_263 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_263 <= REG_262; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_264 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_264 <= REG_263; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_265 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_265 <= REG_264; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_266 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_266 <= REG_265; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_267 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_267 <= REG_266; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_268 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_268 <= REG_267; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_269 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_269 <= REG_268; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_270 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_270 <= REG_269; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_271 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_271 <= REG_270; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_272 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_272 <= REG_271; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_273 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_273 <= REG_272; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_274 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_274 <= REG_273; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_275 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_275 <= REG_274; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_276 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_276 <= REG_275; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_277 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_277 <= REG_276; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_278 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_278 <= REG_277; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_279 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_279 <= REG_278; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_280 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_280 <= REG_279; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_281 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_281 <= REG_280; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_282 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_282 <= REG_281; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_283 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_283 <= REG_282; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_284 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_284 <= REG_283; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_285 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_285 <= REG_284; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_286 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_286 <= REG_285; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_287 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_287 <= REG_286; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_288 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_288 <= REG_287; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_289 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_289 <= REG_288; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_290 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_290 <= REG_289; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_291 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_291 <= REG_290; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_292 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_292 <= REG_291; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_293 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_293 <= REG_292; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_294 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_294 <= REG_293; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_295 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_295 <= REG_294; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_296 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_296 <= REG_295; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_297 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_297 <= REG_296; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_298 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_298 <= REG_297; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_299 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_299 <= REG_298; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_300 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_300 <= REG_299; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_301 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_301 <= REG_300; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_302 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_302 <= REG_301; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_303 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_303 <= REG_302; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_304 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_304 <= REG_303; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_305 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_305 <= REG_304; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_306 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_306 <= REG_305; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_307 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_307 <= REG_306; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_308 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_308 <= REG_307; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_309 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_309 <= REG_308; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_310 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_310 <= REG_309; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_311 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_311 <= REG_310; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_312 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_312 <= REG_311; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_313 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_313 <= REG_312; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_314 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_314 <= REG_313; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_315 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_315 <= REG_314; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_316 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_316 <= REG_315; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_317 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_317 <= REG_316; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_318 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_318 <= REG_317; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_319 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_319 <= REG_318; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_320 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_320 <= REG_319; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_321 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_321 <= REG_320; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_322 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_322 <= REG_321; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_323 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_323 <= REG_322; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_324 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_324 <= REG_323; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_325 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_325 <= REG_324; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_326 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_326 <= REG_325; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_327 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_327 <= REG_326; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_328 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_328 <= REG_327; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_329 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_329 <= REG_328; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_330 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_330 <= REG_329; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_331 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_331 <= REG_330; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_332 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_332 <= REG_331; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_333 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_333 <= REG_332; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_334 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_334 <= REG_333; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_335 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_335 <= REG_334; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_336 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_336 <= REG_335; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_337 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_337 <= REG_336; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_338 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_338 <= REG_337; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_339 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_339 <= REG_338; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_340 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_340 <= REG_339; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_341 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_341 <= REG_340; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_342 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_342 <= REG_341; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_343 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_343 <= REG_342; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_344 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_344 <= REG_343; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_345 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_345 <= REG_344; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_346 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_346 <= REG_345; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_347 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_347 <= REG_346; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_348 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_348 <= REG_347; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_349 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_349 <= REG_348; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_350 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_350 <= REG_349; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_351 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_351 <= REG_350; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_352 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_352 <= REG_351; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_353 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_353 <= REG_352; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_354 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_354 <= REG_353; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_355 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_355 <= REG_354; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_356 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_356 <= REG_355; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_357 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_357 <= REG_356; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_358 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_358 <= REG_357; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_359 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_359 <= REG_358; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_360 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_360 <= REG_359; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_361 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_361 <= REG_360; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_362 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_362 <= REG_361; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_363 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_363 <= REG_362; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_364 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_364 <= REG_363; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_365 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_365 <= REG_364; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_366 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_366 <= REG_365; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_367 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_367 <= REG_366; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_368 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_368 <= REG_367; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_369 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_369 <= REG_368; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_370 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_370 <= REG_369; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_371 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_371 <= REG_370; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_372 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_372 <= REG_371; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_373 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_373 <= REG_372; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_374 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_374 <= REG_373; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_375 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_375 <= REG_374; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_376 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_376 <= REG_375; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_377 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_377 <= REG_376; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_378 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_378 <= REG_377; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_379 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_379 <= REG_378; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_380 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_380 <= REG_379; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_381 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_381 <= REG_380; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_382 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_382 <= REG_381; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_383 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_383 <= REG_382; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_384 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_384 <= REG_383; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_385 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_385 <= REG_384; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_386 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_386 <= REG_385; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_387 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_387 <= REG_386; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_388 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_388 <= REG_387; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_389 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_389 <= REG_388; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_390 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_390 <= REG_389; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_391 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_391 <= REG_390; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_392 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_392 <= REG_391; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_393 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_393 <= REG_392; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_394 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_394 <= REG_393; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_395 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_395 <= REG_394; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_396 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_396 <= REG_395; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_397 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_397 <= REG_396; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_398 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_398 <= REG_397; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_399 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_399 <= REG_398; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_400 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_400 <= REG_399; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_401 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_401 <= REG_400; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_402 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_402 <= REG_401; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_403 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_403 <= REG_402; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_404 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_404 <= REG_403; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_405 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_405 <= REG_404; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_406 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_406 <= REG_405; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_407 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_407 <= REG_406; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_408 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_408 <= REG_407; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_409 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_409 <= REG_408; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_410 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_410 <= REG_409; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_411 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_411 <= REG_410; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_412 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_412 <= REG_411; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_413 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_413 <= REG_412; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_414 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_414 <= REG_413; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_415 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_415 <= REG_414; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_416 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_416 <= REG_415; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_417 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_417 <= REG_416; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_418 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_418 <= REG_417; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_419 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_419 <= REG_418; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_420 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_420 <= REG_419; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_421 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_421 <= REG_420; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_422 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_422 <= REG_421; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_423 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_423 <= REG_422; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_424 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_424 <= REG_423; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_425 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_425 <= REG_424; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_426 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_426 <= REG_425; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_427 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_427 <= REG_426; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_428 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_428 <= REG_427; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_429 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_429 <= REG_428; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_430 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_430 <= REG_429; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_431 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_431 <= REG_430; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_432 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_432 <= REG_431; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_433 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_433 <= REG_432; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_434 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_434 <= REG_433; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_435 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_435 <= REG_434; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_436 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_436 <= REG_435; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_437 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_437 <= REG_436; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_438 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_438 <= REG_437; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_439 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_439 <= REG_438; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_440 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_440 <= REG_439; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_441 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_441 <= REG_440; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_442 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_442 <= REG_441; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_443 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_443 <= REG_442; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_444 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_444 <= REG_443; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_445 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_445 <= REG_444; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_446 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_446 <= REG_445; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_447 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_447 <= REG_446; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_448 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_448 <= REG_447; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_449 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_449 <= REG_448; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_450 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_450 <= REG_449; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_451 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_451 <= REG_450; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_452 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_452 <= REG_451; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_453 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_453 <= REG_452; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_454 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_454 <= REG_453; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_455 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_455 <= REG_454; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_456 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_456 <= REG_455; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_457 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_457 <= REG_456; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_458 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_458 <= REG_457; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_459 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_459 <= REG_458; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_460 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_460 <= REG_459; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_461 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_461 <= REG_460; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_462 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_462 <= REG_461; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_463 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_463 <= REG_462; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_464 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_464 <= REG_463; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_465 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_465 <= REG_464; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_466 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_466 <= REG_465; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_467 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_467 <= REG_466; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_468 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_468 <= REG_467; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_469 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_469 <= REG_468; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_470 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_470 <= REG_469; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_471 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_471 <= REG_470; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_472 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_472 <= REG_471; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_473 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_473 <= REG_472; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_474 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_474 <= REG_473; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_475 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_475 <= REG_474; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_476 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_476 <= REG_475; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_477 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_477 <= REG_476; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_478 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_478 <= REG_477; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_479 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_479 <= REG_478; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_480 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_480 <= REG_479; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_481 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_481 <= REG_480; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_482 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_482 <= REG_481; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_483 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_483 <= REG_482; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_484 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_484 <= REG_483; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_485 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_485 <= REG_484; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_486 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_486 <= REG_485; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_487 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_487 <= REG_486; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_488 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_488 <= REG_487; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_489 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_489 <= REG_488; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_490 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_490 <= REG_489; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_491 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_491 <= REG_490; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_492 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_492 <= REG_491; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_493 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_493 <= REG_492; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_494 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_494 <= REG_493; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_495 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_495 <= REG_494; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_496 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_496 <= REG_495; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_497 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_497 <= REG_496; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_498 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_498 <= REG_497; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_499 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_499 <= REG_498; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_500 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_500 <= REG_499; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_501 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_501 <= REG_500; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_502 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_502 <= REG_501; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_503 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_503 <= REG_502; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_504 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_504 <= REG_503; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_505 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_505 <= REG_504; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_506 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_506 <= REG_505; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_507 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_507 <= REG_506; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_508 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_508 <= REG_507; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_509 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_509 <= REG_508; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_510 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_510 <= REG_509; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_511 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_511 <= REG_510; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_512 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_512 <= REG_511; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_513 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_513 <= REG_512; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_514 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_514 <= REG_513; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_515 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_515 <= REG_514; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_516 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_516 <= REG_515; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_517 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_517 <= REG_516; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_518 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_518 <= REG_517; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_519 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_519 <= REG_518; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_520 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_520 <= REG_519; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_521 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_521 <= REG_520; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_522 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_522 <= REG_521; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_523 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_523 <= REG_522; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_524 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_524 <= REG_523; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_525 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_525 <= REG_524; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_526 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_526 <= REG_525; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_527 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_527 <= REG_526; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_528 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_528 <= REG_527; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_529 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_529 <= REG_528; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_530 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_530 <= REG_529; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_531 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_531 <= REG_530; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_532 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_532 <= REG_531; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_533 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_533 <= REG_532; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_534 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_534 <= REG_533; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_535 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_535 <= REG_534; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_536 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_536 <= REG_535; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_537 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_537 <= REG_536; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_538 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_538 <= REG_537; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_539 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_539 <= REG_538; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_540 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_540 <= REG_539; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_541 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_541 <= REG_540; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_542 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_542 <= REG_541; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_543 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_543 <= REG_542; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_544 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_544 <= REG_543; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_545 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_545 <= REG_544; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_546 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_546 <= REG_545; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_547 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_547 <= REG_546; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_548 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_548 <= REG_547; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_549 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_549 <= REG_548; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_550 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_550 <= REG_549; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_551 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_551 <= REG_550; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_552 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_552 <= REG_551; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_553 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_553 <= REG_552; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_554 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_554 <= REG_553; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_555 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_555 <= REG_554; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_556 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_556 <= REG_555; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_557 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_557 <= REG_556; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_558 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_558 <= REG_557; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_559 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_559 <= REG_558; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_560 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_560 <= REG_559; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_561 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_561 <= REG_560; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_562 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_562 <= REG_561; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_563 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_563 <= REG_562; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_564 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_564 <= REG_563; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_565 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_565 <= REG_564; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_566 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_566 <= REG_565; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_567 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_567 <= REG_566; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_568 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_568 <= REG_567; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_569 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_569 <= REG_568; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_570 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_570 <= REG_569; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_571 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_571 <= REG_570; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_572 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_572 <= REG_571; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_573 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_573 <= REG_572; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_574 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_574 <= REG_573; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_575 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_575 <= REG_574; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_576 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_576 <= REG_575; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_577 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_577 <= REG_576; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_578 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_578 <= REG_577; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_579 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_579 <= REG_578; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_580 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_580 <= REG_579; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_581 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_581 <= REG_580; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_582 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_582 <= REG_581; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_583 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_583 <= REG_582; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_584 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_584 <= REG_583; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_585 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_585 <= REG_584; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_586 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_586 <= REG_585; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_587 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_587 <= REG_586; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_588 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_588 <= REG_587; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_589 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_589 <= REG_588; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_590 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_590 <= REG_589; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_591 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_591 <= REG_590; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_592 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_592 <= REG_591; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_593 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_593 <= REG_592; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_594 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_594 <= REG_593; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_595 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_595 <= REG_594; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_596 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_596 <= REG_595; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_597 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_597 <= REG_596; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_598 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_598 <= REG_597; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_599 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_599 <= REG_598; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_600 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_600 <= REG_599; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_601 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_601 <= REG_600; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_602 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_602 <= REG_601; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_603 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_603 <= REG_602; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_604 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_604 <= REG_603; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_605 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_605 <= REG_604; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_606 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_606 <= REG_605; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_607 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_607 <= REG_606; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_608 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_608 <= REG_607; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_609 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_609 <= REG_608; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_610 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_610 <= REG_609; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_611 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_611 <= REG_610; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_612 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_612 <= REG_611; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_613 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_613 <= REG_612; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_614 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_614 <= REG_613; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_615 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_615 <= REG_614; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_616 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_616 <= REG_615; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_617 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_617 <= REG_616; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_618 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_618 <= REG_617; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_619 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_619 <= REG_618; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_620 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_620 <= REG_619; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_621 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_621 <= REG_620; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_622 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_622 <= REG_621; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_623 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_623 <= REG_622; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_624 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_624 <= REG_623; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_625 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_625 <= REG_624; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_626 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_626 <= REG_625; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_627 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_627 <= REG_626; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_628 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_628 <= REG_627; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_629 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_629 <= REG_628; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_630 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_630 <= REG_629; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_631 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_631 <= REG_630; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_632 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_632 <= REG_631; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_633 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_633 <= REG_632; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_634 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_634 <= REG_633; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_635 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_635 <= REG_634; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_636 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_636 <= REG_635; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_637 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_637 <= REG_636; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_638 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_638 <= REG_637; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_639 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_639 <= REG_638; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_640 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_640 <= REG_639; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_641 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_641 <= REG_640; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_642 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_642 <= REG_641; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_643 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_643 <= REG_642; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_644 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_644 <= REG_643; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_645 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_645 <= REG_644; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_646 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_646 <= REG_645; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_647 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_647 <= REG_646; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_648 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_648 <= REG_647; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_649 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_649 <= REG_648; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_650 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_650 <= REG_649; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_651 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_651 <= REG_650; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_652 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_652 <= REG_651; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_653 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_653 <= REG_652; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_654 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_654 <= REG_653; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_655 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_655 <= REG_654; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_656 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_656 <= REG_655; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_657 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_657 <= REG_656; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_658 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_658 <= REG_657; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_659 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_659 <= REG_658; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_660 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_660 <= REG_659; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_661 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_661 <= REG_660; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_662 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_662 <= REG_661; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_663 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_663 <= REG_662; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_664 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_664 <= REG_663; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_665 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_665 <= REG_664; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_666 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_666 <= REG_665; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_667 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_667 <= REG_666; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_668 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_668 <= REG_667; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_669 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_669 <= REG_668; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_670 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_670 <= REG_669; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_671 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_671 <= REG_670; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_672 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_672 <= REG_671; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_673 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_673 <= REG_672; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_674 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_674 <= REG_673; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_675 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_675 <= REG_674; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_676 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_676 <= REG_675; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_677 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_677 <= REG_676; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_678 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_678 <= REG_677; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_679 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_679 <= REG_678; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_680 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_680 <= REG_679; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_681 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_681 <= REG_680; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_682 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_682 <= REG_681; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_683 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_683 <= REG_682; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_684 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_684 <= REG_683; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_685 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_685 <= REG_684; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_686 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_686 <= REG_685; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_687 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_687 <= REG_686; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_688 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_688 <= REG_687; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_689 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_689 <= REG_688; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_690 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_690 <= REG_689; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_691 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_691 <= REG_690; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_692 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_692 <= REG_691; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_693 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_693 <= REG_692; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_694 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_694 <= REG_693; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_695 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_695 <= REG_694; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_696 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_696 <= REG_695; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_697 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_697 <= REG_696; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_698 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_698 <= REG_697; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_699 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_699 <= REG_698; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_700 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_700 <= REG_699; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_701 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_701 <= REG_700; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_702 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_702 <= REG_701; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_703 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_703 <= REG_702; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_704 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_704 <= REG_703; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_705 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_705 <= REG_704; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_706 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_706 <= REG_705; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_707 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_707 <= REG_706; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_708 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_708 <= REG_707; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_709 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_709 <= REG_708; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_710 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_710 <= REG_709; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_711 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_711 <= REG_710; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_712 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_712 <= REG_711; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_713 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_713 <= REG_712; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_714 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_714 <= REG_713; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_715 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_715 <= REG_714; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_716 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_716 <= REG_715; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_717 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_717 <= REG_716; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_718 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_718 <= REG_717; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_719 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_719 <= REG_718; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_720 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_720 <= REG_719; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_721 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_721 <= REG_720; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_722 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_722 <= REG_721; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_723 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_723 <= REG_722; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_724 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_724 <= REG_723; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_725 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_725 <= REG_724; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_726 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_726 <= REG_725; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_727 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_727 <= REG_726; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_728 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_728 <= REG_727; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_729 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_729 <= REG_728; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_730 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_730 <= REG_729; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_731 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_731 <= REG_730; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_732 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_732 <= REG_731; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_733 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_733 <= REG_732; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_734 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_734 <= REG_733; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_735 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_735 <= REG_734; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_736 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_736 <= REG_735; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_737 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_737 <= REG_736; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_738 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_738 <= REG_737; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_739 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_739 <= REG_738; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_740 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_740 <= REG_739; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_741 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_741 <= REG_740; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_742 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_742 <= REG_741; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_743 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_743 <= REG_742; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_744 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_744 <= REG_743; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_745 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_745 <= REG_744; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_746 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_746 <= REG_745; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_747 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_747 <= REG_746; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_748 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_748 <= REG_747; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_749 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_749 <= REG_748; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_750 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_750 <= REG_749; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_751 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_751 <= REG_750; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_752 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_752 <= REG_751; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_753 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_753 <= REG_752; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_754 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_754 <= REG_753; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_755 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_755 <= REG_754; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_756 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_756 <= REG_755; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_757 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_757 <= REG_756; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_758 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_758 <= REG_757; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_759 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_759 <= REG_758; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_760 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_760 <= REG_759; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_761 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_761 <= REG_760; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_762 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_762 <= REG_761; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_763 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_763 <= REG_762; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_764 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_764 <= REG_763; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_765 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_765 <= REG_764; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_766 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_766 <= REG_765; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_767 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_767 <= REG_766; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_768 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_768 <= REG_767; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_769 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_769 <= REG_768; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_770 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_770 <= REG_769; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_771 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_771 <= REG_770; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_772 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_772 <= REG_771; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_773 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_773 <= REG_772; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_774 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_774 <= REG_773; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_775 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_775 <= REG_774; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_776 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_776 <= REG_775; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_777 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_777 <= REG_776; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_778 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_778 <= REG_777; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_779 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_779 <= REG_778; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_780 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_780 <= REG_779; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_781 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_781 <= REG_780; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_782 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_782 <= REG_781; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_783 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_783 <= REG_782; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_784 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_784 <= REG_783; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_785 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_785 <= REG_784; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_786 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_786 <= REG_785; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_787 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_787 <= REG_786; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_788 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_788 <= REG_787; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_789 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_789 <= REG_788; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_790 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_790 <= REG_789; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_791 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_791 <= REG_790; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_792 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_792 <= REG_791; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_793 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_793 <= REG_792; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_794 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_794 <= REG_793; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_795 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_795 <= REG_794; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_796 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_796 <= REG_795; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_797 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_797 <= REG_796; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_798 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_798 <= REG_797; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_799 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_799 <= REG_798; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_800 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_800 <= REG_799; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_801 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_801 <= REG_800; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_802 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_802 <= REG_801; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_803 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_803 <= REG_802; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_804 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_804 <= REG_803; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_805 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_805 <= REG_804; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_806 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_806 <= REG_805; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_807 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_807 <= REG_806; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_808 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_808 <= REG_807; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_809 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_809 <= REG_808; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_810 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_810 <= REG_809; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_811 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_811 <= REG_810; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_812 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_812 <= REG_811; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_813 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_813 <= REG_812; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_814 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_814 <= REG_813; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_815 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_815 <= REG_814; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_816 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_816 <= REG_815; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_817 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_817 <= REG_816; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_818 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_818 <= REG_817; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_819 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_819 <= REG_818; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_820 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_820 <= REG_819; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_821 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_821 <= REG_820; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_822 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_822 <= REG_821; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_823 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_823 <= REG_822; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_824 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_824 <= REG_823; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_825 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_825 <= REG_824; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_826 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_826 <= REG_825; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_827 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_827 <= REG_826; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_828 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_828 <= REG_827; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_829 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_829 <= REG_828; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_830 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_830 <= REG_829; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_831 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_831 <= REG_830; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_832 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_832 <= REG_831; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_833 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_833 <= REG_832; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_834 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_834 <= REG_833; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_835 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_835 <= REG_834; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_836 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_836 <= REG_835; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_837 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_837 <= REG_836; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_838 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_838 <= REG_837; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_839 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_839 <= REG_838; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_840 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_840 <= REG_839; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_841 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_841 <= REG_840; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_842 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_842 <= REG_841; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_843 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_843 <= REG_842; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_844 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_844 <= REG_843; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_845 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_845 <= REG_844; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_846 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_846 <= REG_845; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_847 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_847 <= REG_846; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_848 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_848 <= REG_847; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_849 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_849 <= REG_848; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_850 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_850 <= REG_849; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_851 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_851 <= REG_850; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_852 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_852 <= REG_851; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_853 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_853 <= REG_852; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_854 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_854 <= REG_853; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_855 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_855 <= REG_854; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_856 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_856 <= REG_855; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_857 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_857 <= REG_856; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_858 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_858 <= REG_857; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_859 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_859 <= REG_858; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_860 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_860 <= REG_859; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_861 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_861 <= REG_860; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_862 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_862 <= REG_861; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_863 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_863 <= REG_862; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_864 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_864 <= REG_863; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_865 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_865 <= REG_864; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_866 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_866 <= REG_865; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_867 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_867 <= REG_866; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_868 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_868 <= REG_867; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_869 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_869 <= REG_868; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_870 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_870 <= REG_869; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_871 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_871 <= REG_870; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_872 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_872 <= REG_871; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_873 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_873 <= REG_872; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_874 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_874 <= REG_873; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_875 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_875 <= REG_874; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_876 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_876 <= REG_875; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_877 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_877 <= REG_876; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_878 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_878 <= REG_877; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_879 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_879 <= REG_878; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_880 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_880 <= REG_879; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_881 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_881 <= REG_880; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_882 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_882 <= REG_881; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_883 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_883 <= REG_882; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_884 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_884 <= REG_883; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_885 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_885 <= REG_884; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_886 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_886 <= REG_885; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_887 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_887 <= REG_886; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_888 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_888 <= REG_887; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_889 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_889 <= REG_888; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_890 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_890 <= REG_889; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_891 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_891 <= REG_890; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_892 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_892 <= REG_891; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_893 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_893 <= REG_892; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_894 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_894 <= REG_893; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_895 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_895 <= REG_894; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_896 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_896 <= REG_895; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_897 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_897 <= REG_896; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_898 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_898 <= REG_897; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_899 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_899 <= REG_898; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_900 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_900 <= REG_899; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_901 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_901 <= REG_900; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_902 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_902 <= REG_901; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_903 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_903 <= REG_902; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_904 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_904 <= REG_903; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_905 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_905 <= REG_904; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_906 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_906 <= REG_905; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_907 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_907 <= REG_906; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_908 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_908 <= REG_907; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_909 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_909 <= REG_908; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_910 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_910 <= REG_909; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_911 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_911 <= REG_910; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_912 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_912 <= REG_911; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_913 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_913 <= REG_912; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_914 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_914 <= REG_913; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_915 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_915 <= REG_914; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_916 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_916 <= REG_915; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_917 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_917 <= REG_916; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_918 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_918 <= REG_917; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_919 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_919 <= REG_918; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_920 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_920 <= REG_919; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_921 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_921 <= REG_920; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_922 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_922 <= REG_921; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_923 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_923 <= REG_922; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_924 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_924 <= REG_923; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_925 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_925 <= REG_924; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_926 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_926 <= REG_925; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_927 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_927 <= REG_926; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_928 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_928 <= REG_927; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_929 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_929 <= REG_928; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_930 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_930 <= REG_929; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_931 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_931 <= REG_930; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_932 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_932 <= REG_931; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_933 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_933 <= REG_932; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_934 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_934 <= REG_933; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_935 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_935 <= REG_934; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_936 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_936 <= REG_935; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_937 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_937 <= REG_936; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_938 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_938 <= REG_937; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_939 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_939 <= REG_938; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_940 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_940 <= REG_939; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_941 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_941 <= REG_940; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_942 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_942 <= REG_941; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_943 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_943 <= REG_942; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_944 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_944 <= REG_943; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_945 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_945 <= REG_944; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_946 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_946 <= REG_945; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_947 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_947 <= REG_946; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_948 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_948 <= REG_947; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_949 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_949 <= REG_948; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_950 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_950 <= REG_949; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_951 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_951 <= REG_950; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_952 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_952 <= REG_951; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_953 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_953 <= REG_952; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_954 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_954 <= REG_953; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_955 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_955 <= REG_954; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_956 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_956 <= REG_955; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_957 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_957 <= REG_956; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_958 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_958 <= REG_957; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_959 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_959 <= REG_958; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_960 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_960 <= REG_959; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_961 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_961 <= REG_960; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_962 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_962 <= REG_961; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_963 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_963 <= REG_962; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_964 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_964 <= REG_963; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_965 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_965 <= REG_964; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_966 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_966 <= REG_965; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_967 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_967 <= REG_966; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_968 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_968 <= REG_967; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_969 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_969 <= REG_968; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_970 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_970 <= REG_969; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_971 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_971 <= REG_970; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_972 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_972 <= REG_971; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_973 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_973 <= REG_972; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_974 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_974 <= REG_973; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_975 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_975 <= REG_974; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_976 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_976 <= REG_975; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_977 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_977 <= REG_976; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_978 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_978 <= REG_977; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_979 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_979 <= REG_978; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_980 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_980 <= REG_979; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_981 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_981 <= REG_980; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_982 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_982 <= REG_981; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_983 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_983 <= REG_982; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_984 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_984 <= REG_983; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_985 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_985 <= REG_984; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_986 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_986 <= REG_985; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_987 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_987 <= REG_986; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_988 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_988 <= REG_987; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_989 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_989 <= REG_988; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_990 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_990 <= REG_989; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_991 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_991 <= REG_990; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_992 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_992 <= REG_991; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_993 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_993 <= REG_992; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_994 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_994 <= REG_993; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_995 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_995 <= REG_994; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_996 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_996 <= REG_995; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_997 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_997 <= REG_996; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      REG_998 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      REG_998 <= REG_997; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[AXI4IntrGenerator.scala 63:23]
      w_fire_1 <= 1'h0; // @[AXI4IntrGenerator.scala 63:23]
    end else begin
      w_fire_1 <= REG_998; // @[AXI4IntrGenerator.scala 63:23]
    end
    if (reset) begin // @[LFSR64.scala 25:23]
      intrGenRegs_6_lfsr <= 64'h1234567887654321; // @[LFSR64.scala 25:23]
    end else if (intrGenRegs_6_lfsr == 64'h0) begin // @[LFSR64.scala 28:18]
      intrGenRegs_6_lfsr <= 64'h1;
    end else begin
      intrGenRegs_6_lfsr <= _intrGenRegs_6_lfsr_T_2;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  value = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  hold_data = _RAND_2[7:0];
  _RAND_3 = {2{`RANDOM}};
  raddr_hold_data = _RAND_3[36:0];
  _RAND_4 = {2{`RANDOM}};
  waddr_hold_data = _RAND_4[36:0];
  _RAND_5 = {1{`RANDOM}};
  bundleIn_0_bid_r = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  bundleIn_0_rid_r = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  intrGenRegs_0 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  intrGenRegs_1 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  intrGenRegs_2 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  intrGenRegs_3 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  intrGenRegs_4 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  intrGenRegs_5 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  intrGenRegs_6 = _RAND_13[31:0];
  _RAND_14 = {2{`RANDOM}};
  randomPosition_lfsr = _RAND_14[63:0];
  _RAND_15 = {1{`RANDOM}};
  REG = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  REG_1 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  REG_2 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  REG_3 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  REG_4 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  REG_5 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  REG_6 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  REG_7 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  REG_8 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  REG_9 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  REG_10 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  REG_11 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  REG_12 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  REG_13 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  REG_14 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  REG_15 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  REG_16 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  REG_17 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  REG_18 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  REG_19 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  REG_20 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  REG_21 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  REG_22 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  REG_23 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  REG_24 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  REG_25 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  REG_26 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  REG_27 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  REG_28 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  REG_29 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  REG_30 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  REG_31 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  REG_32 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  REG_33 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  REG_34 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  REG_35 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  REG_36 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  REG_37 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  REG_38 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  REG_39 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  REG_40 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  REG_41 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  REG_42 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  REG_43 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  REG_44 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  REG_45 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  REG_46 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  REG_47 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  REG_48 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  REG_49 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  REG_50 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  REG_51 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  REG_52 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  REG_53 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  REG_54 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  REG_55 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  REG_56 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  REG_57 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  REG_58 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  REG_59 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  REG_60 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  REG_61 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  REG_62 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  REG_63 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  REG_64 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  REG_65 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  REG_66 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  REG_67 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  REG_68 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  REG_69 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  REG_70 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  REG_71 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  REG_72 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  REG_73 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  REG_74 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  REG_75 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  REG_76 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  REG_77 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  REG_78 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  REG_79 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  REG_80 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  REG_81 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  REG_82 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  REG_83 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  REG_84 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  REG_85 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  REG_86 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  REG_87 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  REG_88 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  REG_89 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  REG_90 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  REG_91 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  REG_92 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  REG_93 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  REG_94 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  REG_95 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  REG_96 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  REG_97 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  REG_98 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  REG_99 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  REG_100 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  REG_101 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  REG_102 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  REG_103 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  REG_104 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  REG_105 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  REG_106 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  REG_107 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  REG_108 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  REG_109 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  REG_110 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  REG_111 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  REG_112 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  REG_113 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  REG_114 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  REG_115 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  REG_116 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  REG_117 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  REG_118 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  REG_119 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  REG_120 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  REG_121 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  REG_122 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  REG_123 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  REG_124 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  REG_125 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  REG_126 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  REG_127 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  REG_128 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  REG_129 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  REG_130 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  REG_131 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  REG_132 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  REG_133 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  REG_134 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  REG_135 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  REG_136 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  REG_137 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  REG_138 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  REG_139 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  REG_140 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  REG_141 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  REG_142 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  REG_143 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  REG_144 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  REG_145 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  REG_146 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  REG_147 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  REG_148 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  REG_149 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  REG_150 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  REG_151 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  REG_152 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  REG_153 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  REG_154 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  REG_155 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  REG_156 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  REG_157 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  REG_158 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  REG_159 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  REG_160 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  REG_161 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  REG_162 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  REG_163 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  REG_164 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  REG_165 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  REG_166 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  REG_167 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  REG_168 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  REG_169 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  REG_170 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  REG_171 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  REG_172 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  REG_173 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  REG_174 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  REG_175 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  REG_176 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  REG_177 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  REG_178 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  REG_179 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  REG_180 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  REG_181 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  REG_182 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  REG_183 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  REG_184 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  REG_185 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  REG_186 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  REG_187 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  REG_188 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  REG_189 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  REG_190 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  REG_191 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  REG_192 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  REG_193 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  REG_194 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  REG_195 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  REG_196 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  REG_197 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  REG_198 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  REG_199 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  REG_200 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  REG_201 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  REG_202 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  REG_203 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  REG_204 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  REG_205 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  REG_206 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  REG_207 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  REG_208 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  REG_209 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  REG_210 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  REG_211 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  REG_212 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  REG_213 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  REG_214 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  REG_215 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  REG_216 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  REG_217 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  REG_218 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  REG_219 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  REG_220 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  REG_221 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  REG_222 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  REG_223 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  REG_224 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  REG_225 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  REG_226 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  REG_227 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  REG_228 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  REG_229 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  REG_230 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  REG_231 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  REG_232 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  REG_233 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  REG_234 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  REG_235 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  REG_236 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  REG_237 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  REG_238 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  REG_239 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  REG_240 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  REG_241 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  REG_242 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  REG_243 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  REG_244 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  REG_245 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  REG_246 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  REG_247 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  REG_248 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  REG_249 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  REG_250 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  REG_251 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  REG_252 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  REG_253 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  REG_254 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  REG_255 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  REG_256 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  REG_257 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  REG_258 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  REG_259 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  REG_260 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  REG_261 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  REG_262 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  REG_263 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  REG_264 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  REG_265 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  REG_266 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  REG_267 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  REG_268 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  REG_269 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  REG_270 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  REG_271 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  REG_272 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  REG_273 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  REG_274 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  REG_275 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  REG_276 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  REG_277 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  REG_278 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  REG_279 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  REG_280 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  REG_281 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  REG_282 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  REG_283 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  REG_284 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  REG_285 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  REG_286 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  REG_287 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  REG_288 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  REG_289 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  REG_290 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  REG_291 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  REG_292 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  REG_293 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  REG_294 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  REG_295 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  REG_296 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  REG_297 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  REG_298 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  REG_299 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  REG_300 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  REG_301 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  REG_302 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  REG_303 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  REG_304 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  REG_305 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  REG_306 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  REG_307 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  REG_308 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  REG_309 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  REG_310 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  REG_311 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  REG_312 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  REG_313 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  REG_314 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  REG_315 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  REG_316 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  REG_317 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  REG_318 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  REG_319 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  REG_320 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  REG_321 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  REG_322 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  REG_323 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  REG_324 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  REG_325 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  REG_326 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  REG_327 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  REG_328 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  REG_329 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  REG_330 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  REG_331 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  REG_332 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  REG_333 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  REG_334 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  REG_335 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  REG_336 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  REG_337 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  REG_338 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  REG_339 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  REG_340 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  REG_341 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  REG_342 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  REG_343 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  REG_344 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  REG_345 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  REG_346 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  REG_347 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  REG_348 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  REG_349 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  REG_350 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  REG_351 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  REG_352 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  REG_353 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  REG_354 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  REG_355 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  REG_356 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  REG_357 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  REG_358 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  REG_359 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  REG_360 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  REG_361 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  REG_362 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  REG_363 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  REG_364 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  REG_365 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  REG_366 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  REG_367 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  REG_368 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  REG_369 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  REG_370 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  REG_371 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  REG_372 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  REG_373 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  REG_374 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  REG_375 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  REG_376 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  REG_377 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  REG_378 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  REG_379 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  REG_380 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  REG_381 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  REG_382 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  REG_383 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  REG_384 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  REG_385 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  REG_386 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  REG_387 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  REG_388 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  REG_389 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  REG_390 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  REG_391 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  REG_392 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  REG_393 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  REG_394 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  REG_395 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  REG_396 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  REG_397 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  REG_398 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  REG_399 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  REG_400 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  REG_401 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  REG_402 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  REG_403 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  REG_404 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  REG_405 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  REG_406 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  REG_407 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  REG_408 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  REG_409 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  REG_410 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  REG_411 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  REG_412 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  REG_413 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  REG_414 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  REG_415 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  REG_416 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  REG_417 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  REG_418 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  REG_419 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  REG_420 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  REG_421 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  REG_422 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  REG_423 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  REG_424 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  REG_425 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  REG_426 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  REG_427 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  REG_428 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  REG_429 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  REG_430 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  REG_431 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  REG_432 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  REG_433 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  REG_434 = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  REG_435 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  REG_436 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  REG_437 = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  REG_438 = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  REG_439 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  REG_440 = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  REG_441 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  REG_442 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  REG_443 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  REG_444 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  REG_445 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  REG_446 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  REG_447 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  REG_448 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  REG_449 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  REG_450 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  REG_451 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  REG_452 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  REG_453 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  REG_454 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  REG_455 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  REG_456 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  REG_457 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  REG_458 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  REG_459 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  REG_460 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  REG_461 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  REG_462 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  REG_463 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  REG_464 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  REG_465 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  REG_466 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  REG_467 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  REG_468 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  REG_469 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  REG_470 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  REG_471 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  REG_472 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  REG_473 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  REG_474 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  REG_475 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  REG_476 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  REG_477 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  REG_478 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  REG_479 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  REG_480 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  REG_481 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  REG_482 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  REG_483 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  REG_484 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  REG_485 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  REG_486 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  REG_487 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  REG_488 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  REG_489 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  REG_490 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  REG_491 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  REG_492 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  REG_493 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  REG_494 = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  REG_495 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  REG_496 = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  REG_497 = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  REG_498 = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  REG_499 = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  REG_500 = _RAND_515[0:0];
  _RAND_516 = {1{`RANDOM}};
  REG_501 = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  REG_502 = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  REG_503 = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  REG_504 = _RAND_519[0:0];
  _RAND_520 = {1{`RANDOM}};
  REG_505 = _RAND_520[0:0];
  _RAND_521 = {1{`RANDOM}};
  REG_506 = _RAND_521[0:0];
  _RAND_522 = {1{`RANDOM}};
  REG_507 = _RAND_522[0:0];
  _RAND_523 = {1{`RANDOM}};
  REG_508 = _RAND_523[0:0];
  _RAND_524 = {1{`RANDOM}};
  REG_509 = _RAND_524[0:0];
  _RAND_525 = {1{`RANDOM}};
  REG_510 = _RAND_525[0:0];
  _RAND_526 = {1{`RANDOM}};
  REG_511 = _RAND_526[0:0];
  _RAND_527 = {1{`RANDOM}};
  REG_512 = _RAND_527[0:0];
  _RAND_528 = {1{`RANDOM}};
  REG_513 = _RAND_528[0:0];
  _RAND_529 = {1{`RANDOM}};
  REG_514 = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  REG_515 = _RAND_530[0:0];
  _RAND_531 = {1{`RANDOM}};
  REG_516 = _RAND_531[0:0];
  _RAND_532 = {1{`RANDOM}};
  REG_517 = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  REG_518 = _RAND_533[0:0];
  _RAND_534 = {1{`RANDOM}};
  REG_519 = _RAND_534[0:0];
  _RAND_535 = {1{`RANDOM}};
  REG_520 = _RAND_535[0:0];
  _RAND_536 = {1{`RANDOM}};
  REG_521 = _RAND_536[0:0];
  _RAND_537 = {1{`RANDOM}};
  REG_522 = _RAND_537[0:0];
  _RAND_538 = {1{`RANDOM}};
  REG_523 = _RAND_538[0:0];
  _RAND_539 = {1{`RANDOM}};
  REG_524 = _RAND_539[0:0];
  _RAND_540 = {1{`RANDOM}};
  REG_525 = _RAND_540[0:0];
  _RAND_541 = {1{`RANDOM}};
  REG_526 = _RAND_541[0:0];
  _RAND_542 = {1{`RANDOM}};
  REG_527 = _RAND_542[0:0];
  _RAND_543 = {1{`RANDOM}};
  REG_528 = _RAND_543[0:0];
  _RAND_544 = {1{`RANDOM}};
  REG_529 = _RAND_544[0:0];
  _RAND_545 = {1{`RANDOM}};
  REG_530 = _RAND_545[0:0];
  _RAND_546 = {1{`RANDOM}};
  REG_531 = _RAND_546[0:0];
  _RAND_547 = {1{`RANDOM}};
  REG_532 = _RAND_547[0:0];
  _RAND_548 = {1{`RANDOM}};
  REG_533 = _RAND_548[0:0];
  _RAND_549 = {1{`RANDOM}};
  REG_534 = _RAND_549[0:0];
  _RAND_550 = {1{`RANDOM}};
  REG_535 = _RAND_550[0:0];
  _RAND_551 = {1{`RANDOM}};
  REG_536 = _RAND_551[0:0];
  _RAND_552 = {1{`RANDOM}};
  REG_537 = _RAND_552[0:0];
  _RAND_553 = {1{`RANDOM}};
  REG_538 = _RAND_553[0:0];
  _RAND_554 = {1{`RANDOM}};
  REG_539 = _RAND_554[0:0];
  _RAND_555 = {1{`RANDOM}};
  REG_540 = _RAND_555[0:0];
  _RAND_556 = {1{`RANDOM}};
  REG_541 = _RAND_556[0:0];
  _RAND_557 = {1{`RANDOM}};
  REG_542 = _RAND_557[0:0];
  _RAND_558 = {1{`RANDOM}};
  REG_543 = _RAND_558[0:0];
  _RAND_559 = {1{`RANDOM}};
  REG_544 = _RAND_559[0:0];
  _RAND_560 = {1{`RANDOM}};
  REG_545 = _RAND_560[0:0];
  _RAND_561 = {1{`RANDOM}};
  REG_546 = _RAND_561[0:0];
  _RAND_562 = {1{`RANDOM}};
  REG_547 = _RAND_562[0:0];
  _RAND_563 = {1{`RANDOM}};
  REG_548 = _RAND_563[0:0];
  _RAND_564 = {1{`RANDOM}};
  REG_549 = _RAND_564[0:0];
  _RAND_565 = {1{`RANDOM}};
  REG_550 = _RAND_565[0:0];
  _RAND_566 = {1{`RANDOM}};
  REG_551 = _RAND_566[0:0];
  _RAND_567 = {1{`RANDOM}};
  REG_552 = _RAND_567[0:0];
  _RAND_568 = {1{`RANDOM}};
  REG_553 = _RAND_568[0:0];
  _RAND_569 = {1{`RANDOM}};
  REG_554 = _RAND_569[0:0];
  _RAND_570 = {1{`RANDOM}};
  REG_555 = _RAND_570[0:0];
  _RAND_571 = {1{`RANDOM}};
  REG_556 = _RAND_571[0:0];
  _RAND_572 = {1{`RANDOM}};
  REG_557 = _RAND_572[0:0];
  _RAND_573 = {1{`RANDOM}};
  REG_558 = _RAND_573[0:0];
  _RAND_574 = {1{`RANDOM}};
  REG_559 = _RAND_574[0:0];
  _RAND_575 = {1{`RANDOM}};
  REG_560 = _RAND_575[0:0];
  _RAND_576 = {1{`RANDOM}};
  REG_561 = _RAND_576[0:0];
  _RAND_577 = {1{`RANDOM}};
  REG_562 = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  REG_563 = _RAND_578[0:0];
  _RAND_579 = {1{`RANDOM}};
  REG_564 = _RAND_579[0:0];
  _RAND_580 = {1{`RANDOM}};
  REG_565 = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  REG_566 = _RAND_581[0:0];
  _RAND_582 = {1{`RANDOM}};
  REG_567 = _RAND_582[0:0];
  _RAND_583 = {1{`RANDOM}};
  REG_568 = _RAND_583[0:0];
  _RAND_584 = {1{`RANDOM}};
  REG_569 = _RAND_584[0:0];
  _RAND_585 = {1{`RANDOM}};
  REG_570 = _RAND_585[0:0];
  _RAND_586 = {1{`RANDOM}};
  REG_571 = _RAND_586[0:0];
  _RAND_587 = {1{`RANDOM}};
  REG_572 = _RAND_587[0:0];
  _RAND_588 = {1{`RANDOM}};
  REG_573 = _RAND_588[0:0];
  _RAND_589 = {1{`RANDOM}};
  REG_574 = _RAND_589[0:0];
  _RAND_590 = {1{`RANDOM}};
  REG_575 = _RAND_590[0:0];
  _RAND_591 = {1{`RANDOM}};
  REG_576 = _RAND_591[0:0];
  _RAND_592 = {1{`RANDOM}};
  REG_577 = _RAND_592[0:0];
  _RAND_593 = {1{`RANDOM}};
  REG_578 = _RAND_593[0:0];
  _RAND_594 = {1{`RANDOM}};
  REG_579 = _RAND_594[0:0];
  _RAND_595 = {1{`RANDOM}};
  REG_580 = _RAND_595[0:0];
  _RAND_596 = {1{`RANDOM}};
  REG_581 = _RAND_596[0:0];
  _RAND_597 = {1{`RANDOM}};
  REG_582 = _RAND_597[0:0];
  _RAND_598 = {1{`RANDOM}};
  REG_583 = _RAND_598[0:0];
  _RAND_599 = {1{`RANDOM}};
  REG_584 = _RAND_599[0:0];
  _RAND_600 = {1{`RANDOM}};
  REG_585 = _RAND_600[0:0];
  _RAND_601 = {1{`RANDOM}};
  REG_586 = _RAND_601[0:0];
  _RAND_602 = {1{`RANDOM}};
  REG_587 = _RAND_602[0:0];
  _RAND_603 = {1{`RANDOM}};
  REG_588 = _RAND_603[0:0];
  _RAND_604 = {1{`RANDOM}};
  REG_589 = _RAND_604[0:0];
  _RAND_605 = {1{`RANDOM}};
  REG_590 = _RAND_605[0:0];
  _RAND_606 = {1{`RANDOM}};
  REG_591 = _RAND_606[0:0];
  _RAND_607 = {1{`RANDOM}};
  REG_592 = _RAND_607[0:0];
  _RAND_608 = {1{`RANDOM}};
  REG_593 = _RAND_608[0:0];
  _RAND_609 = {1{`RANDOM}};
  REG_594 = _RAND_609[0:0];
  _RAND_610 = {1{`RANDOM}};
  REG_595 = _RAND_610[0:0];
  _RAND_611 = {1{`RANDOM}};
  REG_596 = _RAND_611[0:0];
  _RAND_612 = {1{`RANDOM}};
  REG_597 = _RAND_612[0:0];
  _RAND_613 = {1{`RANDOM}};
  REG_598 = _RAND_613[0:0];
  _RAND_614 = {1{`RANDOM}};
  REG_599 = _RAND_614[0:0];
  _RAND_615 = {1{`RANDOM}};
  REG_600 = _RAND_615[0:0];
  _RAND_616 = {1{`RANDOM}};
  REG_601 = _RAND_616[0:0];
  _RAND_617 = {1{`RANDOM}};
  REG_602 = _RAND_617[0:0];
  _RAND_618 = {1{`RANDOM}};
  REG_603 = _RAND_618[0:0];
  _RAND_619 = {1{`RANDOM}};
  REG_604 = _RAND_619[0:0];
  _RAND_620 = {1{`RANDOM}};
  REG_605 = _RAND_620[0:0];
  _RAND_621 = {1{`RANDOM}};
  REG_606 = _RAND_621[0:0];
  _RAND_622 = {1{`RANDOM}};
  REG_607 = _RAND_622[0:0];
  _RAND_623 = {1{`RANDOM}};
  REG_608 = _RAND_623[0:0];
  _RAND_624 = {1{`RANDOM}};
  REG_609 = _RAND_624[0:0];
  _RAND_625 = {1{`RANDOM}};
  REG_610 = _RAND_625[0:0];
  _RAND_626 = {1{`RANDOM}};
  REG_611 = _RAND_626[0:0];
  _RAND_627 = {1{`RANDOM}};
  REG_612 = _RAND_627[0:0];
  _RAND_628 = {1{`RANDOM}};
  REG_613 = _RAND_628[0:0];
  _RAND_629 = {1{`RANDOM}};
  REG_614 = _RAND_629[0:0];
  _RAND_630 = {1{`RANDOM}};
  REG_615 = _RAND_630[0:0];
  _RAND_631 = {1{`RANDOM}};
  REG_616 = _RAND_631[0:0];
  _RAND_632 = {1{`RANDOM}};
  REG_617 = _RAND_632[0:0];
  _RAND_633 = {1{`RANDOM}};
  REG_618 = _RAND_633[0:0];
  _RAND_634 = {1{`RANDOM}};
  REG_619 = _RAND_634[0:0];
  _RAND_635 = {1{`RANDOM}};
  REG_620 = _RAND_635[0:0];
  _RAND_636 = {1{`RANDOM}};
  REG_621 = _RAND_636[0:0];
  _RAND_637 = {1{`RANDOM}};
  REG_622 = _RAND_637[0:0];
  _RAND_638 = {1{`RANDOM}};
  REG_623 = _RAND_638[0:0];
  _RAND_639 = {1{`RANDOM}};
  REG_624 = _RAND_639[0:0];
  _RAND_640 = {1{`RANDOM}};
  REG_625 = _RAND_640[0:0];
  _RAND_641 = {1{`RANDOM}};
  REG_626 = _RAND_641[0:0];
  _RAND_642 = {1{`RANDOM}};
  REG_627 = _RAND_642[0:0];
  _RAND_643 = {1{`RANDOM}};
  REG_628 = _RAND_643[0:0];
  _RAND_644 = {1{`RANDOM}};
  REG_629 = _RAND_644[0:0];
  _RAND_645 = {1{`RANDOM}};
  REG_630 = _RAND_645[0:0];
  _RAND_646 = {1{`RANDOM}};
  REG_631 = _RAND_646[0:0];
  _RAND_647 = {1{`RANDOM}};
  REG_632 = _RAND_647[0:0];
  _RAND_648 = {1{`RANDOM}};
  REG_633 = _RAND_648[0:0];
  _RAND_649 = {1{`RANDOM}};
  REG_634 = _RAND_649[0:0];
  _RAND_650 = {1{`RANDOM}};
  REG_635 = _RAND_650[0:0];
  _RAND_651 = {1{`RANDOM}};
  REG_636 = _RAND_651[0:0];
  _RAND_652 = {1{`RANDOM}};
  REG_637 = _RAND_652[0:0];
  _RAND_653 = {1{`RANDOM}};
  REG_638 = _RAND_653[0:0];
  _RAND_654 = {1{`RANDOM}};
  REG_639 = _RAND_654[0:0];
  _RAND_655 = {1{`RANDOM}};
  REG_640 = _RAND_655[0:0];
  _RAND_656 = {1{`RANDOM}};
  REG_641 = _RAND_656[0:0];
  _RAND_657 = {1{`RANDOM}};
  REG_642 = _RAND_657[0:0];
  _RAND_658 = {1{`RANDOM}};
  REG_643 = _RAND_658[0:0];
  _RAND_659 = {1{`RANDOM}};
  REG_644 = _RAND_659[0:0];
  _RAND_660 = {1{`RANDOM}};
  REG_645 = _RAND_660[0:0];
  _RAND_661 = {1{`RANDOM}};
  REG_646 = _RAND_661[0:0];
  _RAND_662 = {1{`RANDOM}};
  REG_647 = _RAND_662[0:0];
  _RAND_663 = {1{`RANDOM}};
  REG_648 = _RAND_663[0:0];
  _RAND_664 = {1{`RANDOM}};
  REG_649 = _RAND_664[0:0];
  _RAND_665 = {1{`RANDOM}};
  REG_650 = _RAND_665[0:0];
  _RAND_666 = {1{`RANDOM}};
  REG_651 = _RAND_666[0:0];
  _RAND_667 = {1{`RANDOM}};
  REG_652 = _RAND_667[0:0];
  _RAND_668 = {1{`RANDOM}};
  REG_653 = _RAND_668[0:0];
  _RAND_669 = {1{`RANDOM}};
  REG_654 = _RAND_669[0:0];
  _RAND_670 = {1{`RANDOM}};
  REG_655 = _RAND_670[0:0];
  _RAND_671 = {1{`RANDOM}};
  REG_656 = _RAND_671[0:0];
  _RAND_672 = {1{`RANDOM}};
  REG_657 = _RAND_672[0:0];
  _RAND_673 = {1{`RANDOM}};
  REG_658 = _RAND_673[0:0];
  _RAND_674 = {1{`RANDOM}};
  REG_659 = _RAND_674[0:0];
  _RAND_675 = {1{`RANDOM}};
  REG_660 = _RAND_675[0:0];
  _RAND_676 = {1{`RANDOM}};
  REG_661 = _RAND_676[0:0];
  _RAND_677 = {1{`RANDOM}};
  REG_662 = _RAND_677[0:0];
  _RAND_678 = {1{`RANDOM}};
  REG_663 = _RAND_678[0:0];
  _RAND_679 = {1{`RANDOM}};
  REG_664 = _RAND_679[0:0];
  _RAND_680 = {1{`RANDOM}};
  REG_665 = _RAND_680[0:0];
  _RAND_681 = {1{`RANDOM}};
  REG_666 = _RAND_681[0:0];
  _RAND_682 = {1{`RANDOM}};
  REG_667 = _RAND_682[0:0];
  _RAND_683 = {1{`RANDOM}};
  REG_668 = _RAND_683[0:0];
  _RAND_684 = {1{`RANDOM}};
  REG_669 = _RAND_684[0:0];
  _RAND_685 = {1{`RANDOM}};
  REG_670 = _RAND_685[0:0];
  _RAND_686 = {1{`RANDOM}};
  REG_671 = _RAND_686[0:0];
  _RAND_687 = {1{`RANDOM}};
  REG_672 = _RAND_687[0:0];
  _RAND_688 = {1{`RANDOM}};
  REG_673 = _RAND_688[0:0];
  _RAND_689 = {1{`RANDOM}};
  REG_674 = _RAND_689[0:0];
  _RAND_690 = {1{`RANDOM}};
  REG_675 = _RAND_690[0:0];
  _RAND_691 = {1{`RANDOM}};
  REG_676 = _RAND_691[0:0];
  _RAND_692 = {1{`RANDOM}};
  REG_677 = _RAND_692[0:0];
  _RAND_693 = {1{`RANDOM}};
  REG_678 = _RAND_693[0:0];
  _RAND_694 = {1{`RANDOM}};
  REG_679 = _RAND_694[0:0];
  _RAND_695 = {1{`RANDOM}};
  REG_680 = _RAND_695[0:0];
  _RAND_696 = {1{`RANDOM}};
  REG_681 = _RAND_696[0:0];
  _RAND_697 = {1{`RANDOM}};
  REG_682 = _RAND_697[0:0];
  _RAND_698 = {1{`RANDOM}};
  REG_683 = _RAND_698[0:0];
  _RAND_699 = {1{`RANDOM}};
  REG_684 = _RAND_699[0:0];
  _RAND_700 = {1{`RANDOM}};
  REG_685 = _RAND_700[0:0];
  _RAND_701 = {1{`RANDOM}};
  REG_686 = _RAND_701[0:0];
  _RAND_702 = {1{`RANDOM}};
  REG_687 = _RAND_702[0:0];
  _RAND_703 = {1{`RANDOM}};
  REG_688 = _RAND_703[0:0];
  _RAND_704 = {1{`RANDOM}};
  REG_689 = _RAND_704[0:0];
  _RAND_705 = {1{`RANDOM}};
  REG_690 = _RAND_705[0:0];
  _RAND_706 = {1{`RANDOM}};
  REG_691 = _RAND_706[0:0];
  _RAND_707 = {1{`RANDOM}};
  REG_692 = _RAND_707[0:0];
  _RAND_708 = {1{`RANDOM}};
  REG_693 = _RAND_708[0:0];
  _RAND_709 = {1{`RANDOM}};
  REG_694 = _RAND_709[0:0];
  _RAND_710 = {1{`RANDOM}};
  REG_695 = _RAND_710[0:0];
  _RAND_711 = {1{`RANDOM}};
  REG_696 = _RAND_711[0:0];
  _RAND_712 = {1{`RANDOM}};
  REG_697 = _RAND_712[0:0];
  _RAND_713 = {1{`RANDOM}};
  REG_698 = _RAND_713[0:0];
  _RAND_714 = {1{`RANDOM}};
  REG_699 = _RAND_714[0:0];
  _RAND_715 = {1{`RANDOM}};
  REG_700 = _RAND_715[0:0];
  _RAND_716 = {1{`RANDOM}};
  REG_701 = _RAND_716[0:0];
  _RAND_717 = {1{`RANDOM}};
  REG_702 = _RAND_717[0:0];
  _RAND_718 = {1{`RANDOM}};
  REG_703 = _RAND_718[0:0];
  _RAND_719 = {1{`RANDOM}};
  REG_704 = _RAND_719[0:0];
  _RAND_720 = {1{`RANDOM}};
  REG_705 = _RAND_720[0:0];
  _RAND_721 = {1{`RANDOM}};
  REG_706 = _RAND_721[0:0];
  _RAND_722 = {1{`RANDOM}};
  REG_707 = _RAND_722[0:0];
  _RAND_723 = {1{`RANDOM}};
  REG_708 = _RAND_723[0:0];
  _RAND_724 = {1{`RANDOM}};
  REG_709 = _RAND_724[0:0];
  _RAND_725 = {1{`RANDOM}};
  REG_710 = _RAND_725[0:0];
  _RAND_726 = {1{`RANDOM}};
  REG_711 = _RAND_726[0:0];
  _RAND_727 = {1{`RANDOM}};
  REG_712 = _RAND_727[0:0];
  _RAND_728 = {1{`RANDOM}};
  REG_713 = _RAND_728[0:0];
  _RAND_729 = {1{`RANDOM}};
  REG_714 = _RAND_729[0:0];
  _RAND_730 = {1{`RANDOM}};
  REG_715 = _RAND_730[0:0];
  _RAND_731 = {1{`RANDOM}};
  REG_716 = _RAND_731[0:0];
  _RAND_732 = {1{`RANDOM}};
  REG_717 = _RAND_732[0:0];
  _RAND_733 = {1{`RANDOM}};
  REG_718 = _RAND_733[0:0];
  _RAND_734 = {1{`RANDOM}};
  REG_719 = _RAND_734[0:0];
  _RAND_735 = {1{`RANDOM}};
  REG_720 = _RAND_735[0:0];
  _RAND_736 = {1{`RANDOM}};
  REG_721 = _RAND_736[0:0];
  _RAND_737 = {1{`RANDOM}};
  REG_722 = _RAND_737[0:0];
  _RAND_738 = {1{`RANDOM}};
  REG_723 = _RAND_738[0:0];
  _RAND_739 = {1{`RANDOM}};
  REG_724 = _RAND_739[0:0];
  _RAND_740 = {1{`RANDOM}};
  REG_725 = _RAND_740[0:0];
  _RAND_741 = {1{`RANDOM}};
  REG_726 = _RAND_741[0:0];
  _RAND_742 = {1{`RANDOM}};
  REG_727 = _RAND_742[0:0];
  _RAND_743 = {1{`RANDOM}};
  REG_728 = _RAND_743[0:0];
  _RAND_744 = {1{`RANDOM}};
  REG_729 = _RAND_744[0:0];
  _RAND_745 = {1{`RANDOM}};
  REG_730 = _RAND_745[0:0];
  _RAND_746 = {1{`RANDOM}};
  REG_731 = _RAND_746[0:0];
  _RAND_747 = {1{`RANDOM}};
  REG_732 = _RAND_747[0:0];
  _RAND_748 = {1{`RANDOM}};
  REG_733 = _RAND_748[0:0];
  _RAND_749 = {1{`RANDOM}};
  REG_734 = _RAND_749[0:0];
  _RAND_750 = {1{`RANDOM}};
  REG_735 = _RAND_750[0:0];
  _RAND_751 = {1{`RANDOM}};
  REG_736 = _RAND_751[0:0];
  _RAND_752 = {1{`RANDOM}};
  REG_737 = _RAND_752[0:0];
  _RAND_753 = {1{`RANDOM}};
  REG_738 = _RAND_753[0:0];
  _RAND_754 = {1{`RANDOM}};
  REG_739 = _RAND_754[0:0];
  _RAND_755 = {1{`RANDOM}};
  REG_740 = _RAND_755[0:0];
  _RAND_756 = {1{`RANDOM}};
  REG_741 = _RAND_756[0:0];
  _RAND_757 = {1{`RANDOM}};
  REG_742 = _RAND_757[0:0];
  _RAND_758 = {1{`RANDOM}};
  REG_743 = _RAND_758[0:0];
  _RAND_759 = {1{`RANDOM}};
  REG_744 = _RAND_759[0:0];
  _RAND_760 = {1{`RANDOM}};
  REG_745 = _RAND_760[0:0];
  _RAND_761 = {1{`RANDOM}};
  REG_746 = _RAND_761[0:0];
  _RAND_762 = {1{`RANDOM}};
  REG_747 = _RAND_762[0:0];
  _RAND_763 = {1{`RANDOM}};
  REG_748 = _RAND_763[0:0];
  _RAND_764 = {1{`RANDOM}};
  REG_749 = _RAND_764[0:0];
  _RAND_765 = {1{`RANDOM}};
  REG_750 = _RAND_765[0:0];
  _RAND_766 = {1{`RANDOM}};
  REG_751 = _RAND_766[0:0];
  _RAND_767 = {1{`RANDOM}};
  REG_752 = _RAND_767[0:0];
  _RAND_768 = {1{`RANDOM}};
  REG_753 = _RAND_768[0:0];
  _RAND_769 = {1{`RANDOM}};
  REG_754 = _RAND_769[0:0];
  _RAND_770 = {1{`RANDOM}};
  REG_755 = _RAND_770[0:0];
  _RAND_771 = {1{`RANDOM}};
  REG_756 = _RAND_771[0:0];
  _RAND_772 = {1{`RANDOM}};
  REG_757 = _RAND_772[0:0];
  _RAND_773 = {1{`RANDOM}};
  REG_758 = _RAND_773[0:0];
  _RAND_774 = {1{`RANDOM}};
  REG_759 = _RAND_774[0:0];
  _RAND_775 = {1{`RANDOM}};
  REG_760 = _RAND_775[0:0];
  _RAND_776 = {1{`RANDOM}};
  REG_761 = _RAND_776[0:0];
  _RAND_777 = {1{`RANDOM}};
  REG_762 = _RAND_777[0:0];
  _RAND_778 = {1{`RANDOM}};
  REG_763 = _RAND_778[0:0];
  _RAND_779 = {1{`RANDOM}};
  REG_764 = _RAND_779[0:0];
  _RAND_780 = {1{`RANDOM}};
  REG_765 = _RAND_780[0:0];
  _RAND_781 = {1{`RANDOM}};
  REG_766 = _RAND_781[0:0];
  _RAND_782 = {1{`RANDOM}};
  REG_767 = _RAND_782[0:0];
  _RAND_783 = {1{`RANDOM}};
  REG_768 = _RAND_783[0:0];
  _RAND_784 = {1{`RANDOM}};
  REG_769 = _RAND_784[0:0];
  _RAND_785 = {1{`RANDOM}};
  REG_770 = _RAND_785[0:0];
  _RAND_786 = {1{`RANDOM}};
  REG_771 = _RAND_786[0:0];
  _RAND_787 = {1{`RANDOM}};
  REG_772 = _RAND_787[0:0];
  _RAND_788 = {1{`RANDOM}};
  REG_773 = _RAND_788[0:0];
  _RAND_789 = {1{`RANDOM}};
  REG_774 = _RAND_789[0:0];
  _RAND_790 = {1{`RANDOM}};
  REG_775 = _RAND_790[0:0];
  _RAND_791 = {1{`RANDOM}};
  REG_776 = _RAND_791[0:0];
  _RAND_792 = {1{`RANDOM}};
  REG_777 = _RAND_792[0:0];
  _RAND_793 = {1{`RANDOM}};
  REG_778 = _RAND_793[0:0];
  _RAND_794 = {1{`RANDOM}};
  REG_779 = _RAND_794[0:0];
  _RAND_795 = {1{`RANDOM}};
  REG_780 = _RAND_795[0:0];
  _RAND_796 = {1{`RANDOM}};
  REG_781 = _RAND_796[0:0];
  _RAND_797 = {1{`RANDOM}};
  REG_782 = _RAND_797[0:0];
  _RAND_798 = {1{`RANDOM}};
  REG_783 = _RAND_798[0:0];
  _RAND_799 = {1{`RANDOM}};
  REG_784 = _RAND_799[0:0];
  _RAND_800 = {1{`RANDOM}};
  REG_785 = _RAND_800[0:0];
  _RAND_801 = {1{`RANDOM}};
  REG_786 = _RAND_801[0:0];
  _RAND_802 = {1{`RANDOM}};
  REG_787 = _RAND_802[0:0];
  _RAND_803 = {1{`RANDOM}};
  REG_788 = _RAND_803[0:0];
  _RAND_804 = {1{`RANDOM}};
  REG_789 = _RAND_804[0:0];
  _RAND_805 = {1{`RANDOM}};
  REG_790 = _RAND_805[0:0];
  _RAND_806 = {1{`RANDOM}};
  REG_791 = _RAND_806[0:0];
  _RAND_807 = {1{`RANDOM}};
  REG_792 = _RAND_807[0:0];
  _RAND_808 = {1{`RANDOM}};
  REG_793 = _RAND_808[0:0];
  _RAND_809 = {1{`RANDOM}};
  REG_794 = _RAND_809[0:0];
  _RAND_810 = {1{`RANDOM}};
  REG_795 = _RAND_810[0:0];
  _RAND_811 = {1{`RANDOM}};
  REG_796 = _RAND_811[0:0];
  _RAND_812 = {1{`RANDOM}};
  REG_797 = _RAND_812[0:0];
  _RAND_813 = {1{`RANDOM}};
  REG_798 = _RAND_813[0:0];
  _RAND_814 = {1{`RANDOM}};
  REG_799 = _RAND_814[0:0];
  _RAND_815 = {1{`RANDOM}};
  REG_800 = _RAND_815[0:0];
  _RAND_816 = {1{`RANDOM}};
  REG_801 = _RAND_816[0:0];
  _RAND_817 = {1{`RANDOM}};
  REG_802 = _RAND_817[0:0];
  _RAND_818 = {1{`RANDOM}};
  REG_803 = _RAND_818[0:0];
  _RAND_819 = {1{`RANDOM}};
  REG_804 = _RAND_819[0:0];
  _RAND_820 = {1{`RANDOM}};
  REG_805 = _RAND_820[0:0];
  _RAND_821 = {1{`RANDOM}};
  REG_806 = _RAND_821[0:0];
  _RAND_822 = {1{`RANDOM}};
  REG_807 = _RAND_822[0:0];
  _RAND_823 = {1{`RANDOM}};
  REG_808 = _RAND_823[0:0];
  _RAND_824 = {1{`RANDOM}};
  REG_809 = _RAND_824[0:0];
  _RAND_825 = {1{`RANDOM}};
  REG_810 = _RAND_825[0:0];
  _RAND_826 = {1{`RANDOM}};
  REG_811 = _RAND_826[0:0];
  _RAND_827 = {1{`RANDOM}};
  REG_812 = _RAND_827[0:0];
  _RAND_828 = {1{`RANDOM}};
  REG_813 = _RAND_828[0:0];
  _RAND_829 = {1{`RANDOM}};
  REG_814 = _RAND_829[0:0];
  _RAND_830 = {1{`RANDOM}};
  REG_815 = _RAND_830[0:0];
  _RAND_831 = {1{`RANDOM}};
  REG_816 = _RAND_831[0:0];
  _RAND_832 = {1{`RANDOM}};
  REG_817 = _RAND_832[0:0];
  _RAND_833 = {1{`RANDOM}};
  REG_818 = _RAND_833[0:0];
  _RAND_834 = {1{`RANDOM}};
  REG_819 = _RAND_834[0:0];
  _RAND_835 = {1{`RANDOM}};
  REG_820 = _RAND_835[0:0];
  _RAND_836 = {1{`RANDOM}};
  REG_821 = _RAND_836[0:0];
  _RAND_837 = {1{`RANDOM}};
  REG_822 = _RAND_837[0:0];
  _RAND_838 = {1{`RANDOM}};
  REG_823 = _RAND_838[0:0];
  _RAND_839 = {1{`RANDOM}};
  REG_824 = _RAND_839[0:0];
  _RAND_840 = {1{`RANDOM}};
  REG_825 = _RAND_840[0:0];
  _RAND_841 = {1{`RANDOM}};
  REG_826 = _RAND_841[0:0];
  _RAND_842 = {1{`RANDOM}};
  REG_827 = _RAND_842[0:0];
  _RAND_843 = {1{`RANDOM}};
  REG_828 = _RAND_843[0:0];
  _RAND_844 = {1{`RANDOM}};
  REG_829 = _RAND_844[0:0];
  _RAND_845 = {1{`RANDOM}};
  REG_830 = _RAND_845[0:0];
  _RAND_846 = {1{`RANDOM}};
  REG_831 = _RAND_846[0:0];
  _RAND_847 = {1{`RANDOM}};
  REG_832 = _RAND_847[0:0];
  _RAND_848 = {1{`RANDOM}};
  REG_833 = _RAND_848[0:0];
  _RAND_849 = {1{`RANDOM}};
  REG_834 = _RAND_849[0:0];
  _RAND_850 = {1{`RANDOM}};
  REG_835 = _RAND_850[0:0];
  _RAND_851 = {1{`RANDOM}};
  REG_836 = _RAND_851[0:0];
  _RAND_852 = {1{`RANDOM}};
  REG_837 = _RAND_852[0:0];
  _RAND_853 = {1{`RANDOM}};
  REG_838 = _RAND_853[0:0];
  _RAND_854 = {1{`RANDOM}};
  REG_839 = _RAND_854[0:0];
  _RAND_855 = {1{`RANDOM}};
  REG_840 = _RAND_855[0:0];
  _RAND_856 = {1{`RANDOM}};
  REG_841 = _RAND_856[0:0];
  _RAND_857 = {1{`RANDOM}};
  REG_842 = _RAND_857[0:0];
  _RAND_858 = {1{`RANDOM}};
  REG_843 = _RAND_858[0:0];
  _RAND_859 = {1{`RANDOM}};
  REG_844 = _RAND_859[0:0];
  _RAND_860 = {1{`RANDOM}};
  REG_845 = _RAND_860[0:0];
  _RAND_861 = {1{`RANDOM}};
  REG_846 = _RAND_861[0:0];
  _RAND_862 = {1{`RANDOM}};
  REG_847 = _RAND_862[0:0];
  _RAND_863 = {1{`RANDOM}};
  REG_848 = _RAND_863[0:0];
  _RAND_864 = {1{`RANDOM}};
  REG_849 = _RAND_864[0:0];
  _RAND_865 = {1{`RANDOM}};
  REG_850 = _RAND_865[0:0];
  _RAND_866 = {1{`RANDOM}};
  REG_851 = _RAND_866[0:0];
  _RAND_867 = {1{`RANDOM}};
  REG_852 = _RAND_867[0:0];
  _RAND_868 = {1{`RANDOM}};
  REG_853 = _RAND_868[0:0];
  _RAND_869 = {1{`RANDOM}};
  REG_854 = _RAND_869[0:0];
  _RAND_870 = {1{`RANDOM}};
  REG_855 = _RAND_870[0:0];
  _RAND_871 = {1{`RANDOM}};
  REG_856 = _RAND_871[0:0];
  _RAND_872 = {1{`RANDOM}};
  REG_857 = _RAND_872[0:0];
  _RAND_873 = {1{`RANDOM}};
  REG_858 = _RAND_873[0:0];
  _RAND_874 = {1{`RANDOM}};
  REG_859 = _RAND_874[0:0];
  _RAND_875 = {1{`RANDOM}};
  REG_860 = _RAND_875[0:0];
  _RAND_876 = {1{`RANDOM}};
  REG_861 = _RAND_876[0:0];
  _RAND_877 = {1{`RANDOM}};
  REG_862 = _RAND_877[0:0];
  _RAND_878 = {1{`RANDOM}};
  REG_863 = _RAND_878[0:0];
  _RAND_879 = {1{`RANDOM}};
  REG_864 = _RAND_879[0:0];
  _RAND_880 = {1{`RANDOM}};
  REG_865 = _RAND_880[0:0];
  _RAND_881 = {1{`RANDOM}};
  REG_866 = _RAND_881[0:0];
  _RAND_882 = {1{`RANDOM}};
  REG_867 = _RAND_882[0:0];
  _RAND_883 = {1{`RANDOM}};
  REG_868 = _RAND_883[0:0];
  _RAND_884 = {1{`RANDOM}};
  REG_869 = _RAND_884[0:0];
  _RAND_885 = {1{`RANDOM}};
  REG_870 = _RAND_885[0:0];
  _RAND_886 = {1{`RANDOM}};
  REG_871 = _RAND_886[0:0];
  _RAND_887 = {1{`RANDOM}};
  REG_872 = _RAND_887[0:0];
  _RAND_888 = {1{`RANDOM}};
  REG_873 = _RAND_888[0:0];
  _RAND_889 = {1{`RANDOM}};
  REG_874 = _RAND_889[0:0];
  _RAND_890 = {1{`RANDOM}};
  REG_875 = _RAND_890[0:0];
  _RAND_891 = {1{`RANDOM}};
  REG_876 = _RAND_891[0:0];
  _RAND_892 = {1{`RANDOM}};
  REG_877 = _RAND_892[0:0];
  _RAND_893 = {1{`RANDOM}};
  REG_878 = _RAND_893[0:0];
  _RAND_894 = {1{`RANDOM}};
  REG_879 = _RAND_894[0:0];
  _RAND_895 = {1{`RANDOM}};
  REG_880 = _RAND_895[0:0];
  _RAND_896 = {1{`RANDOM}};
  REG_881 = _RAND_896[0:0];
  _RAND_897 = {1{`RANDOM}};
  REG_882 = _RAND_897[0:0];
  _RAND_898 = {1{`RANDOM}};
  REG_883 = _RAND_898[0:0];
  _RAND_899 = {1{`RANDOM}};
  REG_884 = _RAND_899[0:0];
  _RAND_900 = {1{`RANDOM}};
  REG_885 = _RAND_900[0:0];
  _RAND_901 = {1{`RANDOM}};
  REG_886 = _RAND_901[0:0];
  _RAND_902 = {1{`RANDOM}};
  REG_887 = _RAND_902[0:0];
  _RAND_903 = {1{`RANDOM}};
  REG_888 = _RAND_903[0:0];
  _RAND_904 = {1{`RANDOM}};
  REG_889 = _RAND_904[0:0];
  _RAND_905 = {1{`RANDOM}};
  REG_890 = _RAND_905[0:0];
  _RAND_906 = {1{`RANDOM}};
  REG_891 = _RAND_906[0:0];
  _RAND_907 = {1{`RANDOM}};
  REG_892 = _RAND_907[0:0];
  _RAND_908 = {1{`RANDOM}};
  REG_893 = _RAND_908[0:0];
  _RAND_909 = {1{`RANDOM}};
  REG_894 = _RAND_909[0:0];
  _RAND_910 = {1{`RANDOM}};
  REG_895 = _RAND_910[0:0];
  _RAND_911 = {1{`RANDOM}};
  REG_896 = _RAND_911[0:0];
  _RAND_912 = {1{`RANDOM}};
  REG_897 = _RAND_912[0:0];
  _RAND_913 = {1{`RANDOM}};
  REG_898 = _RAND_913[0:0];
  _RAND_914 = {1{`RANDOM}};
  REG_899 = _RAND_914[0:0];
  _RAND_915 = {1{`RANDOM}};
  REG_900 = _RAND_915[0:0];
  _RAND_916 = {1{`RANDOM}};
  REG_901 = _RAND_916[0:0];
  _RAND_917 = {1{`RANDOM}};
  REG_902 = _RAND_917[0:0];
  _RAND_918 = {1{`RANDOM}};
  REG_903 = _RAND_918[0:0];
  _RAND_919 = {1{`RANDOM}};
  REG_904 = _RAND_919[0:0];
  _RAND_920 = {1{`RANDOM}};
  REG_905 = _RAND_920[0:0];
  _RAND_921 = {1{`RANDOM}};
  REG_906 = _RAND_921[0:0];
  _RAND_922 = {1{`RANDOM}};
  REG_907 = _RAND_922[0:0];
  _RAND_923 = {1{`RANDOM}};
  REG_908 = _RAND_923[0:0];
  _RAND_924 = {1{`RANDOM}};
  REG_909 = _RAND_924[0:0];
  _RAND_925 = {1{`RANDOM}};
  REG_910 = _RAND_925[0:0];
  _RAND_926 = {1{`RANDOM}};
  REG_911 = _RAND_926[0:0];
  _RAND_927 = {1{`RANDOM}};
  REG_912 = _RAND_927[0:0];
  _RAND_928 = {1{`RANDOM}};
  REG_913 = _RAND_928[0:0];
  _RAND_929 = {1{`RANDOM}};
  REG_914 = _RAND_929[0:0];
  _RAND_930 = {1{`RANDOM}};
  REG_915 = _RAND_930[0:0];
  _RAND_931 = {1{`RANDOM}};
  REG_916 = _RAND_931[0:0];
  _RAND_932 = {1{`RANDOM}};
  REG_917 = _RAND_932[0:0];
  _RAND_933 = {1{`RANDOM}};
  REG_918 = _RAND_933[0:0];
  _RAND_934 = {1{`RANDOM}};
  REG_919 = _RAND_934[0:0];
  _RAND_935 = {1{`RANDOM}};
  REG_920 = _RAND_935[0:0];
  _RAND_936 = {1{`RANDOM}};
  REG_921 = _RAND_936[0:0];
  _RAND_937 = {1{`RANDOM}};
  REG_922 = _RAND_937[0:0];
  _RAND_938 = {1{`RANDOM}};
  REG_923 = _RAND_938[0:0];
  _RAND_939 = {1{`RANDOM}};
  REG_924 = _RAND_939[0:0];
  _RAND_940 = {1{`RANDOM}};
  REG_925 = _RAND_940[0:0];
  _RAND_941 = {1{`RANDOM}};
  REG_926 = _RAND_941[0:0];
  _RAND_942 = {1{`RANDOM}};
  REG_927 = _RAND_942[0:0];
  _RAND_943 = {1{`RANDOM}};
  REG_928 = _RAND_943[0:0];
  _RAND_944 = {1{`RANDOM}};
  REG_929 = _RAND_944[0:0];
  _RAND_945 = {1{`RANDOM}};
  REG_930 = _RAND_945[0:0];
  _RAND_946 = {1{`RANDOM}};
  REG_931 = _RAND_946[0:0];
  _RAND_947 = {1{`RANDOM}};
  REG_932 = _RAND_947[0:0];
  _RAND_948 = {1{`RANDOM}};
  REG_933 = _RAND_948[0:0];
  _RAND_949 = {1{`RANDOM}};
  REG_934 = _RAND_949[0:0];
  _RAND_950 = {1{`RANDOM}};
  REG_935 = _RAND_950[0:0];
  _RAND_951 = {1{`RANDOM}};
  REG_936 = _RAND_951[0:0];
  _RAND_952 = {1{`RANDOM}};
  REG_937 = _RAND_952[0:0];
  _RAND_953 = {1{`RANDOM}};
  REG_938 = _RAND_953[0:0];
  _RAND_954 = {1{`RANDOM}};
  REG_939 = _RAND_954[0:0];
  _RAND_955 = {1{`RANDOM}};
  REG_940 = _RAND_955[0:0];
  _RAND_956 = {1{`RANDOM}};
  REG_941 = _RAND_956[0:0];
  _RAND_957 = {1{`RANDOM}};
  REG_942 = _RAND_957[0:0];
  _RAND_958 = {1{`RANDOM}};
  REG_943 = _RAND_958[0:0];
  _RAND_959 = {1{`RANDOM}};
  REG_944 = _RAND_959[0:0];
  _RAND_960 = {1{`RANDOM}};
  REG_945 = _RAND_960[0:0];
  _RAND_961 = {1{`RANDOM}};
  REG_946 = _RAND_961[0:0];
  _RAND_962 = {1{`RANDOM}};
  REG_947 = _RAND_962[0:0];
  _RAND_963 = {1{`RANDOM}};
  REG_948 = _RAND_963[0:0];
  _RAND_964 = {1{`RANDOM}};
  REG_949 = _RAND_964[0:0];
  _RAND_965 = {1{`RANDOM}};
  REG_950 = _RAND_965[0:0];
  _RAND_966 = {1{`RANDOM}};
  REG_951 = _RAND_966[0:0];
  _RAND_967 = {1{`RANDOM}};
  REG_952 = _RAND_967[0:0];
  _RAND_968 = {1{`RANDOM}};
  REG_953 = _RAND_968[0:0];
  _RAND_969 = {1{`RANDOM}};
  REG_954 = _RAND_969[0:0];
  _RAND_970 = {1{`RANDOM}};
  REG_955 = _RAND_970[0:0];
  _RAND_971 = {1{`RANDOM}};
  REG_956 = _RAND_971[0:0];
  _RAND_972 = {1{`RANDOM}};
  REG_957 = _RAND_972[0:0];
  _RAND_973 = {1{`RANDOM}};
  REG_958 = _RAND_973[0:0];
  _RAND_974 = {1{`RANDOM}};
  REG_959 = _RAND_974[0:0];
  _RAND_975 = {1{`RANDOM}};
  REG_960 = _RAND_975[0:0];
  _RAND_976 = {1{`RANDOM}};
  REG_961 = _RAND_976[0:0];
  _RAND_977 = {1{`RANDOM}};
  REG_962 = _RAND_977[0:0];
  _RAND_978 = {1{`RANDOM}};
  REG_963 = _RAND_978[0:0];
  _RAND_979 = {1{`RANDOM}};
  REG_964 = _RAND_979[0:0];
  _RAND_980 = {1{`RANDOM}};
  REG_965 = _RAND_980[0:0];
  _RAND_981 = {1{`RANDOM}};
  REG_966 = _RAND_981[0:0];
  _RAND_982 = {1{`RANDOM}};
  REG_967 = _RAND_982[0:0];
  _RAND_983 = {1{`RANDOM}};
  REG_968 = _RAND_983[0:0];
  _RAND_984 = {1{`RANDOM}};
  REG_969 = _RAND_984[0:0];
  _RAND_985 = {1{`RANDOM}};
  REG_970 = _RAND_985[0:0];
  _RAND_986 = {1{`RANDOM}};
  REG_971 = _RAND_986[0:0];
  _RAND_987 = {1{`RANDOM}};
  REG_972 = _RAND_987[0:0];
  _RAND_988 = {1{`RANDOM}};
  REG_973 = _RAND_988[0:0];
  _RAND_989 = {1{`RANDOM}};
  REG_974 = _RAND_989[0:0];
  _RAND_990 = {1{`RANDOM}};
  REG_975 = _RAND_990[0:0];
  _RAND_991 = {1{`RANDOM}};
  REG_976 = _RAND_991[0:0];
  _RAND_992 = {1{`RANDOM}};
  REG_977 = _RAND_992[0:0];
  _RAND_993 = {1{`RANDOM}};
  REG_978 = _RAND_993[0:0];
  _RAND_994 = {1{`RANDOM}};
  REG_979 = _RAND_994[0:0];
  _RAND_995 = {1{`RANDOM}};
  REG_980 = _RAND_995[0:0];
  _RAND_996 = {1{`RANDOM}};
  REG_981 = _RAND_996[0:0];
  _RAND_997 = {1{`RANDOM}};
  REG_982 = _RAND_997[0:0];
  _RAND_998 = {1{`RANDOM}};
  REG_983 = _RAND_998[0:0];
  _RAND_999 = {1{`RANDOM}};
  REG_984 = _RAND_999[0:0];
  _RAND_1000 = {1{`RANDOM}};
  REG_985 = _RAND_1000[0:0];
  _RAND_1001 = {1{`RANDOM}};
  REG_986 = _RAND_1001[0:0];
  _RAND_1002 = {1{`RANDOM}};
  REG_987 = _RAND_1002[0:0];
  _RAND_1003 = {1{`RANDOM}};
  REG_988 = _RAND_1003[0:0];
  _RAND_1004 = {1{`RANDOM}};
  REG_989 = _RAND_1004[0:0];
  _RAND_1005 = {1{`RANDOM}};
  REG_990 = _RAND_1005[0:0];
  _RAND_1006 = {1{`RANDOM}};
  REG_991 = _RAND_1006[0:0];
  _RAND_1007 = {1{`RANDOM}};
  REG_992 = _RAND_1007[0:0];
  _RAND_1008 = {1{`RANDOM}};
  REG_993 = _RAND_1008[0:0];
  _RAND_1009 = {1{`RANDOM}};
  REG_994 = _RAND_1009[0:0];
  _RAND_1010 = {1{`RANDOM}};
  REG_995 = _RAND_1010[0:0];
  _RAND_1011 = {1{`RANDOM}};
  REG_996 = _RAND_1011[0:0];
  _RAND_1012 = {1{`RANDOM}};
  REG_997 = _RAND_1012[0:0];
  _RAND_1013 = {1{`RANDOM}};
  REG_998 = _RAND_1013[0:0];
  _RAND_1014 = {1{`RANDOM}};
  w_fire_1 = _RAND_1014[0:0];
  _RAND_1015 = {2{`RANDOM}};
  intrGenRegs_6_lfsr = _RAND_1015[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

