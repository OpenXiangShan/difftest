/***************************************************************************************
* Copyright (c) 2025 Beijing Institute of Open Source Chip (BOSC)
* Copyright (c) 2020-2025 Institute of Computing Technology, Chinese Academy of Sciences
*
* DiffTest is licensed under Mulan PSL v2.
* You can use this software according to the terms and conditions of the Mulan PSL v2.
* You may obtain a copy of Mulan PSL v2 at:
*          http://license.coscl.org.cn/MulanPSL2
*
* THIS SOFTWARE IS PROVIDED ON AN "AS IS" BASIS, WITHOUT WARRANTIES OF ANY KIND,
* EITHER EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO NON-INFRINGEMENT,
* MERCHANTABILITY OR FIT FOR A PARTICULAR PURPOSE.
*
* See the Mulan PSL v2 for more details.
***************************************************************************************/

module DifftestClockGate(
	input     CK,
	input	    E,
	output    Q
);

`ifdef SYNTHESIS
	BUFGCE bufgce_1 (
		.O(Q),
		.I(CK),
		.CE(E)
	);
`else
	reg EN;
	always_latch begin
		if (!CK) EN = E;
	end
	assign Q = CK & EN;
`endif // SYNTHESIS
endmodule
