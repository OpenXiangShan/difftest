module DelayN_36(
  input         clock,
  input  [31:0] io_in,
  output [31:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] REG; // @[Hold.scala 89:18]
  reg [31:0] REG_1; // @[Hold.scala 89:18]
  reg [31:0] REG_2; // @[Hold.scala 89:18]
  reg [31:0] REG_3; // @[Hold.scala 89:18]
  reg [31:0] REG_4; // @[Hold.scala 89:18]
  reg [31:0] REG_5; // @[Hold.scala 89:18]
  reg [31:0] REG_6; // @[Hold.scala 89:18]
  reg [31:0] REG_7; // @[Hold.scala 89:18]
  reg [31:0] REG_8; // @[Hold.scala 89:18]
  reg [31:0] REG_9; // @[Hold.scala 89:18]
  reg [31:0] REG_10; // @[Hold.scala 89:18]
  reg [31:0] REG_11; // @[Hold.scala 89:18]
  reg [31:0] REG_12; // @[Hold.scala 89:18]
  reg [31:0] REG_13; // @[Hold.scala 89:18]
  reg [31:0] REG_14; // @[Hold.scala 89:18]
  reg [31:0] REG_15; // @[Hold.scala 89:18]
  reg [31:0] REG_16; // @[Hold.scala 89:18]
  reg [31:0] REG_17; // @[Hold.scala 89:18]
  reg [31:0] REG_18; // @[Hold.scala 89:18]
  reg [31:0] REG_19; // @[Hold.scala 89:18]
  reg [31:0] REG_20; // @[Hold.scala 89:18]
  reg [31:0] REG_21; // @[Hold.scala 89:18]
  reg [31:0] REG_22; // @[Hold.scala 89:18]
  reg [31:0] REG_23; // @[Hold.scala 89:18]
  reg [31:0] REG_24; // @[Hold.scala 89:18]
  reg [31:0] REG_25; // @[Hold.scala 89:18]
  reg [31:0] REG_26; // @[Hold.scala 89:18]
  reg [31:0] REG_27; // @[Hold.scala 89:18]
  reg [31:0] REG_28; // @[Hold.scala 89:18]
  reg [31:0] REG_29; // @[Hold.scala 89:18]
  reg [31:0] REG_30; // @[Hold.scala 89:18]
  reg [31:0] REG_31; // @[Hold.scala 89:18]
  reg [31:0] REG_32; // @[Hold.scala 89:18]
  reg [31:0] REG_33; // @[Hold.scala 89:18]
  reg [31:0] REG_34; // @[Hold.scala 89:18]
  reg [31:0] REG_35; // @[Hold.scala 89:18]
  reg [31:0] REG_36; // @[Hold.scala 89:18]
  reg [31:0] REG_37; // @[Hold.scala 89:18]
  reg [31:0] REG_38; // @[Hold.scala 89:18]
  reg [31:0] REG_39; // @[Hold.scala 89:18]
  reg [31:0] REG_40; // @[Hold.scala 89:18]
  reg [31:0] REG_41; // @[Hold.scala 89:18]
  reg [31:0] REG_42; // @[Hold.scala 89:18]
  reg [31:0] REG_43; // @[Hold.scala 89:18]
  reg [31:0] REG_44; // @[Hold.scala 89:18]
  reg [31:0] REG_45; // @[Hold.scala 89:18]
  reg [31:0] REG_46; // @[Hold.scala 89:18]
  reg [31:0] REG_47; // @[Hold.scala 89:18]
  reg [31:0] REG_48; // @[Hold.scala 89:18]
  reg [31:0] REG_49; // @[Hold.scala 89:18]
  reg [31:0] REG_50; // @[Hold.scala 89:18]
  reg [31:0] REG_51; // @[Hold.scala 89:18]
  reg [31:0] REG_52; // @[Hold.scala 89:18]
  reg [31:0] REG_53; // @[Hold.scala 89:18]
  reg [31:0] REG_54; // @[Hold.scala 89:18]
  reg [31:0] REG_55; // @[Hold.scala 89:18]
  reg [31:0] REG_56; // @[Hold.scala 89:18]
  reg [31:0] REG_57; // @[Hold.scala 89:18]
  reg [31:0] REG_58; // @[Hold.scala 89:18]
  reg [31:0] REG_59; // @[Hold.scala 89:18]
  reg [31:0] REG_60; // @[Hold.scala 89:18]
  reg [31:0] REG_61; // @[Hold.scala 89:18]
  reg [31:0] REG_62; // @[Hold.scala 89:18]
  reg [31:0] REG_63; // @[Hold.scala 89:18]
  reg [31:0] REG_64; // @[Hold.scala 89:18]
  reg [31:0] REG_65; // @[Hold.scala 89:18]
  reg [31:0] REG_66; // @[Hold.scala 89:18]
  reg [31:0] REG_67; // @[Hold.scala 89:18]
  reg [31:0] REG_68; // @[Hold.scala 89:18]
  reg [31:0] REG_69; // @[Hold.scala 89:18]
  reg [31:0] REG_70; // @[Hold.scala 89:18]
  reg [31:0] REG_71; // @[Hold.scala 89:18]
  reg [31:0] REG_72; // @[Hold.scala 89:18]
  reg [31:0] REG_73; // @[Hold.scala 89:18]
  reg [31:0] REG_74; // @[Hold.scala 89:18]
  reg [31:0] REG_75; // @[Hold.scala 89:18]
  reg [31:0] REG_76; // @[Hold.scala 89:18]
  reg [31:0] REG_77; // @[Hold.scala 89:18]
  reg [31:0] REG_78; // @[Hold.scala 89:18]
  reg [31:0] REG_79; // @[Hold.scala 89:18]
  reg [31:0] REG_80; // @[Hold.scala 89:18]
  reg [31:0] REG_81; // @[Hold.scala 89:18]
  reg [31:0] REG_82; // @[Hold.scala 89:18]
  reg [31:0] REG_83; // @[Hold.scala 89:18]
  reg [31:0] REG_84; // @[Hold.scala 89:18]
  reg [31:0] REG_85; // @[Hold.scala 89:18]
  reg [31:0] REG_86; // @[Hold.scala 89:18]
  reg [31:0] REG_87; // @[Hold.scala 89:18]
  reg [31:0] REG_88; // @[Hold.scala 89:18]
  reg [31:0] REG_89; // @[Hold.scala 89:18]
  reg [31:0] REG_90; // @[Hold.scala 89:18]
  reg [31:0] REG_91; // @[Hold.scala 89:18]
  reg [31:0] REG_92; // @[Hold.scala 89:18]
  reg [31:0] REG_93; // @[Hold.scala 89:18]
  reg [31:0] REG_94; // @[Hold.scala 89:18]
  reg [31:0] REG_95; // @[Hold.scala 89:18]
  reg [31:0] REG_96; // @[Hold.scala 89:18]
  reg [31:0] REG_97; // @[Hold.scala 89:18]
  reg [31:0] REG_98; // @[Hold.scala 89:18]
  reg [31:0] REG_99; // @[Hold.scala 89:18]
  reg [31:0] REG_100; // @[Hold.scala 89:18]
  reg [31:0] REG_101; // @[Hold.scala 89:18]
  reg [31:0] REG_102; // @[Hold.scala 89:18]
  reg [31:0] REG_103; // @[Hold.scala 89:18]
  reg [31:0] REG_104; // @[Hold.scala 89:18]
  reg [31:0] REG_105; // @[Hold.scala 89:18]
  reg [31:0] REG_106; // @[Hold.scala 89:18]
  reg [31:0] REG_107; // @[Hold.scala 89:18]
  reg [31:0] REG_108; // @[Hold.scala 89:18]
  reg [31:0] REG_109; // @[Hold.scala 89:18]
  reg [31:0] REG_110; // @[Hold.scala 89:18]
  reg [31:0] REG_111; // @[Hold.scala 89:18]
  reg [31:0] REG_112; // @[Hold.scala 89:18]
  reg [31:0] REG_113; // @[Hold.scala 89:18]
  reg [31:0] REG_114; // @[Hold.scala 89:18]
  reg [31:0] REG_115; // @[Hold.scala 89:18]
  reg [31:0] REG_116; // @[Hold.scala 89:18]
  reg [31:0] REG_117; // @[Hold.scala 89:18]
  reg [31:0] REG_118; // @[Hold.scala 89:18]
  reg [31:0] REG_119; // @[Hold.scala 89:18]
  reg [31:0] REG_120; // @[Hold.scala 89:18]
  reg [31:0] REG_121; // @[Hold.scala 89:18]
  reg [31:0] REG_122; // @[Hold.scala 89:18]
  reg [31:0] REG_123; // @[Hold.scala 89:18]
  reg [31:0] REG_124; // @[Hold.scala 89:18]
  reg [31:0] REG_125; // @[Hold.scala 89:18]
  reg [31:0] REG_126; // @[Hold.scala 89:18]
  reg [31:0] REG_127; // @[Hold.scala 89:18]
  reg [31:0] REG_128; // @[Hold.scala 89:18]
  reg [31:0] REG_129; // @[Hold.scala 89:18]
  reg [31:0] REG_130; // @[Hold.scala 89:18]
  reg [31:0] REG_131; // @[Hold.scala 89:18]
  reg [31:0] REG_132; // @[Hold.scala 89:18]
  reg [31:0] REG_133; // @[Hold.scala 89:18]
  reg [31:0] REG_134; // @[Hold.scala 89:18]
  reg [31:0] REG_135; // @[Hold.scala 89:18]
  reg [31:0] REG_136; // @[Hold.scala 89:18]
  reg [31:0] REG_137; // @[Hold.scala 89:18]
  reg [31:0] REG_138; // @[Hold.scala 89:18]
  reg [31:0] REG_139; // @[Hold.scala 89:18]
  reg [31:0] REG_140; // @[Hold.scala 89:18]
  reg [31:0] REG_141; // @[Hold.scala 89:18]
  reg [31:0] REG_142; // @[Hold.scala 89:18]
  reg [31:0] REG_143; // @[Hold.scala 89:18]
  reg [31:0] REG_144; // @[Hold.scala 89:18]
  reg [31:0] REG_145; // @[Hold.scala 89:18]
  reg [31:0] REG_146; // @[Hold.scala 89:18]
  reg [31:0] REG_147; // @[Hold.scala 89:18]
  reg [31:0] REG_148; // @[Hold.scala 89:18]
  reg [31:0] REG_149; // @[Hold.scala 89:18]
  reg [31:0] REG_150; // @[Hold.scala 89:18]
  reg [31:0] REG_151; // @[Hold.scala 89:18]
  reg [31:0] REG_152; // @[Hold.scala 89:18]
  reg [31:0] REG_153; // @[Hold.scala 89:18]
  reg [31:0] REG_154; // @[Hold.scala 89:18]
  reg [31:0] REG_155; // @[Hold.scala 89:18]
  reg [31:0] REG_156; // @[Hold.scala 89:18]
  reg [31:0] REG_157; // @[Hold.scala 89:18]
  reg [31:0] REG_158; // @[Hold.scala 89:18]
  reg [31:0] REG_159; // @[Hold.scala 89:18]
  reg [31:0] REG_160; // @[Hold.scala 89:18]
  reg [31:0] REG_161; // @[Hold.scala 89:18]
  reg [31:0] REG_162; // @[Hold.scala 89:18]
  reg [31:0] REG_163; // @[Hold.scala 89:18]
  reg [31:0] REG_164; // @[Hold.scala 89:18]
  reg [31:0] REG_165; // @[Hold.scala 89:18]
  reg [31:0] REG_166; // @[Hold.scala 89:18]
  reg [31:0] REG_167; // @[Hold.scala 89:18]
  reg [31:0] REG_168; // @[Hold.scala 89:18]
  reg [31:0] REG_169; // @[Hold.scala 89:18]
  reg [31:0] REG_170; // @[Hold.scala 89:18]
  reg [31:0] REG_171; // @[Hold.scala 89:18]
  reg [31:0] REG_172; // @[Hold.scala 89:18]
  reg [31:0] REG_173; // @[Hold.scala 89:18]
  reg [31:0] REG_174; // @[Hold.scala 89:18]
  reg [31:0] REG_175; // @[Hold.scala 89:18]
  reg [31:0] REG_176; // @[Hold.scala 89:18]
  reg [31:0] REG_177; // @[Hold.scala 89:18]
  reg [31:0] REG_178; // @[Hold.scala 89:18]
  reg [31:0] REG_179; // @[Hold.scala 89:18]
  reg [31:0] REG_180; // @[Hold.scala 89:18]
  reg [31:0] REG_181; // @[Hold.scala 89:18]
  reg [31:0] REG_182; // @[Hold.scala 89:18]
  reg [31:0] REG_183; // @[Hold.scala 89:18]
  reg [31:0] REG_184; // @[Hold.scala 89:18]
  reg [31:0] REG_185; // @[Hold.scala 89:18]
  reg [31:0] REG_186; // @[Hold.scala 89:18]
  reg [31:0] REG_187; // @[Hold.scala 89:18]
  reg [31:0] REG_188; // @[Hold.scala 89:18]
  reg [31:0] REG_189; // @[Hold.scala 89:18]
  reg [31:0] REG_190; // @[Hold.scala 89:18]
  reg [31:0] REG_191; // @[Hold.scala 89:18]
  reg [31:0] REG_192; // @[Hold.scala 89:18]
  reg [31:0] REG_193; // @[Hold.scala 89:18]
  reg [31:0] REG_194; // @[Hold.scala 89:18]
  reg [31:0] REG_195; // @[Hold.scala 89:18]
  reg [31:0] REG_196; // @[Hold.scala 89:18]
  reg [31:0] REG_197; // @[Hold.scala 89:18]
  reg [31:0] REG_198; // @[Hold.scala 89:18]
  reg [31:0] REG_199; // @[Hold.scala 89:18]
  reg [31:0] REG_200; // @[Hold.scala 89:18]
  reg [31:0] REG_201; // @[Hold.scala 89:18]
  reg [31:0] REG_202; // @[Hold.scala 89:18]
  reg [31:0] REG_203; // @[Hold.scala 89:18]
  reg [31:0] REG_204; // @[Hold.scala 89:18]
  reg [31:0] REG_205; // @[Hold.scala 89:18]
  reg [31:0] REG_206; // @[Hold.scala 89:18]
  reg [31:0] REG_207; // @[Hold.scala 89:18]
  reg [31:0] REG_208; // @[Hold.scala 89:18]
  reg [31:0] REG_209; // @[Hold.scala 89:18]
  reg [31:0] REG_210; // @[Hold.scala 89:18]
  reg [31:0] REG_211; // @[Hold.scala 89:18]
  reg [31:0] REG_212; // @[Hold.scala 89:18]
  reg [31:0] REG_213; // @[Hold.scala 89:18]
  reg [31:0] REG_214; // @[Hold.scala 89:18]
  reg [31:0] REG_215; // @[Hold.scala 89:18]
  reg [31:0] REG_216; // @[Hold.scala 89:18]
  reg [31:0] REG_217; // @[Hold.scala 89:18]
  reg [31:0] REG_218; // @[Hold.scala 89:18]
  reg [31:0] REG_219; // @[Hold.scala 89:18]
  reg [31:0] REG_220; // @[Hold.scala 89:18]
  reg [31:0] REG_221; // @[Hold.scala 89:18]
  reg [31:0] REG_222; // @[Hold.scala 89:18]
  reg [31:0] REG_223; // @[Hold.scala 89:18]
  reg [31:0] REG_224; // @[Hold.scala 89:18]
  reg [31:0] REG_225; // @[Hold.scala 89:18]
  reg [31:0] REG_226; // @[Hold.scala 89:18]
  reg [31:0] REG_227; // @[Hold.scala 89:18]
  reg [31:0] REG_228; // @[Hold.scala 89:18]
  reg [31:0] REG_229; // @[Hold.scala 89:18]
  reg [31:0] REG_230; // @[Hold.scala 89:18]
  reg [31:0] REG_231; // @[Hold.scala 89:18]
  reg [31:0] REG_232; // @[Hold.scala 89:18]
  reg [31:0] REG_233; // @[Hold.scala 89:18]
  reg [31:0] REG_234; // @[Hold.scala 89:18]
  reg [31:0] REG_235; // @[Hold.scala 89:18]
  reg [31:0] REG_236; // @[Hold.scala 89:18]
  reg [31:0] REG_237; // @[Hold.scala 89:18]
  reg [31:0] REG_238; // @[Hold.scala 89:18]
  reg [31:0] REG_239; // @[Hold.scala 89:18]
  reg [31:0] REG_240; // @[Hold.scala 89:18]
  reg [31:0] REG_241; // @[Hold.scala 89:18]
  reg [31:0] REG_242; // @[Hold.scala 89:18]
  reg [31:0] REG_243; // @[Hold.scala 89:18]
  reg [31:0] REG_244; // @[Hold.scala 89:18]
  reg [31:0] REG_245; // @[Hold.scala 89:18]
  reg [31:0] REG_246; // @[Hold.scala 89:18]
  reg [31:0] REG_247; // @[Hold.scala 89:18]
  reg [31:0] REG_248; // @[Hold.scala 89:18]
  reg [31:0] REG_249; // @[Hold.scala 89:18]
  reg [31:0] REG_250; // @[Hold.scala 89:18]
  reg [31:0] REG_251; // @[Hold.scala 89:18]
  reg [31:0] REG_252; // @[Hold.scala 89:18]
  reg [31:0] REG_253; // @[Hold.scala 89:18]
  reg [31:0] REG_254; // @[Hold.scala 89:18]
  reg [31:0] REG_255; // @[Hold.scala 89:18]
  reg [31:0] REG_256; // @[Hold.scala 89:18]
  reg [31:0] REG_257; // @[Hold.scala 89:18]
  reg [31:0] REG_258; // @[Hold.scala 89:18]
  reg [31:0] REG_259; // @[Hold.scala 89:18]
  reg [31:0] REG_260; // @[Hold.scala 89:18]
  reg [31:0] REG_261; // @[Hold.scala 89:18]
  reg [31:0] REG_262; // @[Hold.scala 89:18]
  reg [31:0] REG_263; // @[Hold.scala 89:18]
  reg [31:0] REG_264; // @[Hold.scala 89:18]
  reg [31:0] REG_265; // @[Hold.scala 89:18]
  reg [31:0] REG_266; // @[Hold.scala 89:18]
  reg [31:0] REG_267; // @[Hold.scala 89:18]
  reg [31:0] REG_268; // @[Hold.scala 89:18]
  reg [31:0] REG_269; // @[Hold.scala 89:18]
  reg [31:0] REG_270; // @[Hold.scala 89:18]
  reg [31:0] REG_271; // @[Hold.scala 89:18]
  reg [31:0] REG_272; // @[Hold.scala 89:18]
  reg [31:0] REG_273; // @[Hold.scala 89:18]
  reg [31:0] REG_274; // @[Hold.scala 89:18]
  reg [31:0] REG_275; // @[Hold.scala 89:18]
  reg [31:0] REG_276; // @[Hold.scala 89:18]
  reg [31:0] REG_277; // @[Hold.scala 89:18]
  reg [31:0] REG_278; // @[Hold.scala 89:18]
  reg [31:0] REG_279; // @[Hold.scala 89:18]
  reg [31:0] REG_280; // @[Hold.scala 89:18]
  reg [31:0] REG_281; // @[Hold.scala 89:18]
  reg [31:0] REG_282; // @[Hold.scala 89:18]
  reg [31:0] REG_283; // @[Hold.scala 89:18]
  reg [31:0] REG_284; // @[Hold.scala 89:18]
  reg [31:0] REG_285; // @[Hold.scala 89:18]
  reg [31:0] REG_286; // @[Hold.scala 89:18]
  reg [31:0] REG_287; // @[Hold.scala 89:18]
  reg [31:0] REG_288; // @[Hold.scala 89:18]
  reg [31:0] REG_289; // @[Hold.scala 89:18]
  reg [31:0] REG_290; // @[Hold.scala 89:18]
  reg [31:0] REG_291; // @[Hold.scala 89:18]
  reg [31:0] REG_292; // @[Hold.scala 89:18]
  reg [31:0] REG_293; // @[Hold.scala 89:18]
  reg [31:0] REG_294; // @[Hold.scala 89:18]
  reg [31:0] REG_295; // @[Hold.scala 89:18]
  reg [31:0] REG_296; // @[Hold.scala 89:18]
  reg [31:0] REG_297; // @[Hold.scala 89:18]
  reg [31:0] REG_298; // @[Hold.scala 89:18]
  reg [31:0] REG_299; // @[Hold.scala 89:18]
  reg [31:0] REG_300; // @[Hold.scala 89:18]
  reg [31:0] REG_301; // @[Hold.scala 89:18]
  reg [31:0] REG_302; // @[Hold.scala 89:18]
  reg [31:0] REG_303; // @[Hold.scala 89:18]
  reg [31:0] REG_304; // @[Hold.scala 89:18]
  reg [31:0] REG_305; // @[Hold.scala 89:18]
  reg [31:0] REG_306; // @[Hold.scala 89:18]
  reg [31:0] REG_307; // @[Hold.scala 89:18]
  reg [31:0] REG_308; // @[Hold.scala 89:18]
  reg [31:0] REG_309; // @[Hold.scala 89:18]
  reg [31:0] REG_310; // @[Hold.scala 89:18]
  reg [31:0] REG_311; // @[Hold.scala 89:18]
  reg [31:0] REG_312; // @[Hold.scala 89:18]
  reg [31:0] REG_313; // @[Hold.scala 89:18]
  reg [31:0] REG_314; // @[Hold.scala 89:18]
  reg [31:0] REG_315; // @[Hold.scala 89:18]
  reg [31:0] REG_316; // @[Hold.scala 89:18]
  reg [31:0] REG_317; // @[Hold.scala 89:18]
  reg [31:0] REG_318; // @[Hold.scala 89:18]
  reg [31:0] REG_319; // @[Hold.scala 89:18]
  reg [31:0] REG_320; // @[Hold.scala 89:18]
  reg [31:0] REG_321; // @[Hold.scala 89:18]
  reg [31:0] REG_322; // @[Hold.scala 89:18]
  reg [31:0] REG_323; // @[Hold.scala 89:18]
  reg [31:0] REG_324; // @[Hold.scala 89:18]
  reg [31:0] REG_325; // @[Hold.scala 89:18]
  reg [31:0] REG_326; // @[Hold.scala 89:18]
  reg [31:0] REG_327; // @[Hold.scala 89:18]
  reg [31:0] REG_328; // @[Hold.scala 89:18]
  reg [31:0] REG_329; // @[Hold.scala 89:18]
  reg [31:0] REG_330; // @[Hold.scala 89:18]
  reg [31:0] REG_331; // @[Hold.scala 89:18]
  reg [31:0] REG_332; // @[Hold.scala 89:18]
  reg [31:0] REG_333; // @[Hold.scala 89:18]
  reg [31:0] REG_334; // @[Hold.scala 89:18]
  reg [31:0] REG_335; // @[Hold.scala 89:18]
  reg [31:0] REG_336; // @[Hold.scala 89:18]
  reg [31:0] REG_337; // @[Hold.scala 89:18]
  reg [31:0] REG_338; // @[Hold.scala 89:18]
  reg [31:0] REG_339; // @[Hold.scala 89:18]
  reg [31:0] REG_340; // @[Hold.scala 89:18]
  reg [31:0] REG_341; // @[Hold.scala 89:18]
  reg [31:0] REG_342; // @[Hold.scala 89:18]
  reg [31:0] REG_343; // @[Hold.scala 89:18]
  reg [31:0] REG_344; // @[Hold.scala 89:18]
  reg [31:0] REG_345; // @[Hold.scala 89:18]
  reg [31:0] REG_346; // @[Hold.scala 89:18]
  reg [31:0] REG_347; // @[Hold.scala 89:18]
  reg [31:0] REG_348; // @[Hold.scala 89:18]
  reg [31:0] REG_349; // @[Hold.scala 89:18]
  reg [31:0] REG_350; // @[Hold.scala 89:18]
  reg [31:0] REG_351; // @[Hold.scala 89:18]
  reg [31:0] REG_352; // @[Hold.scala 89:18]
  reg [31:0] REG_353; // @[Hold.scala 89:18]
  reg [31:0] REG_354; // @[Hold.scala 89:18]
  reg [31:0] REG_355; // @[Hold.scala 89:18]
  reg [31:0] REG_356; // @[Hold.scala 89:18]
  reg [31:0] REG_357; // @[Hold.scala 89:18]
  reg [31:0] REG_358; // @[Hold.scala 89:18]
  reg [31:0] REG_359; // @[Hold.scala 89:18]
  reg [31:0] REG_360; // @[Hold.scala 89:18]
  reg [31:0] REG_361; // @[Hold.scala 89:18]
  reg [31:0] REG_362; // @[Hold.scala 89:18]
  reg [31:0] REG_363; // @[Hold.scala 89:18]
  reg [31:0] REG_364; // @[Hold.scala 89:18]
  reg [31:0] REG_365; // @[Hold.scala 89:18]
  reg [31:0] REG_366; // @[Hold.scala 89:18]
  reg [31:0] REG_367; // @[Hold.scala 89:18]
  reg [31:0] REG_368; // @[Hold.scala 89:18]
  reg [31:0] REG_369; // @[Hold.scala 89:18]
  reg [31:0] REG_370; // @[Hold.scala 89:18]
  reg [31:0] REG_371; // @[Hold.scala 89:18]
  reg [31:0] REG_372; // @[Hold.scala 89:18]
  reg [31:0] REG_373; // @[Hold.scala 89:18]
  reg [31:0] REG_374; // @[Hold.scala 89:18]
  reg [31:0] REG_375; // @[Hold.scala 89:18]
  reg [31:0] REG_376; // @[Hold.scala 89:18]
  reg [31:0] REG_377; // @[Hold.scala 89:18]
  reg [31:0] REG_378; // @[Hold.scala 89:18]
  reg [31:0] REG_379; // @[Hold.scala 89:18]
  reg [31:0] REG_380; // @[Hold.scala 89:18]
  reg [31:0] REG_381; // @[Hold.scala 89:18]
  reg [31:0] REG_382; // @[Hold.scala 89:18]
  reg [31:0] REG_383; // @[Hold.scala 89:18]
  reg [31:0] REG_384; // @[Hold.scala 89:18]
  reg [31:0] REG_385; // @[Hold.scala 89:18]
  reg [31:0] REG_386; // @[Hold.scala 89:18]
  reg [31:0] REG_387; // @[Hold.scala 89:18]
  reg [31:0] REG_388; // @[Hold.scala 89:18]
  reg [31:0] REG_389; // @[Hold.scala 89:18]
  reg [31:0] REG_390; // @[Hold.scala 89:18]
  reg [31:0] REG_391; // @[Hold.scala 89:18]
  reg [31:0] REG_392; // @[Hold.scala 89:18]
  reg [31:0] REG_393; // @[Hold.scala 89:18]
  reg [31:0] REG_394; // @[Hold.scala 89:18]
  reg [31:0] REG_395; // @[Hold.scala 89:18]
  reg [31:0] REG_396; // @[Hold.scala 89:18]
  reg [31:0] REG_397; // @[Hold.scala 89:18]
  reg [31:0] REG_398; // @[Hold.scala 89:18]
  reg [31:0] REG_399; // @[Hold.scala 89:18]
  reg [31:0] REG_400; // @[Hold.scala 89:18]
  reg [31:0] REG_401; // @[Hold.scala 89:18]
  reg [31:0] REG_402; // @[Hold.scala 89:18]
  reg [31:0] REG_403; // @[Hold.scala 89:18]
  reg [31:0] REG_404; // @[Hold.scala 89:18]
  reg [31:0] REG_405; // @[Hold.scala 89:18]
  reg [31:0] REG_406; // @[Hold.scala 89:18]
  reg [31:0] REG_407; // @[Hold.scala 89:18]
  reg [31:0] REG_408; // @[Hold.scala 89:18]
  reg [31:0] REG_409; // @[Hold.scala 89:18]
  reg [31:0] REG_410; // @[Hold.scala 89:18]
  reg [31:0] REG_411; // @[Hold.scala 89:18]
  reg [31:0] REG_412; // @[Hold.scala 89:18]
  reg [31:0] REG_413; // @[Hold.scala 89:18]
  reg [31:0] REG_414; // @[Hold.scala 89:18]
  reg [31:0] REG_415; // @[Hold.scala 89:18]
  reg [31:0] REG_416; // @[Hold.scala 89:18]
  reg [31:0] REG_417; // @[Hold.scala 89:18]
  reg [31:0] REG_418; // @[Hold.scala 89:18]
  reg [31:0] REG_419; // @[Hold.scala 89:18]
  reg [31:0] REG_420; // @[Hold.scala 89:18]
  reg [31:0] REG_421; // @[Hold.scala 89:18]
  reg [31:0] REG_422; // @[Hold.scala 89:18]
  reg [31:0] REG_423; // @[Hold.scala 89:18]
  reg [31:0] REG_424; // @[Hold.scala 89:18]
  reg [31:0] REG_425; // @[Hold.scala 89:18]
  reg [31:0] REG_426; // @[Hold.scala 89:18]
  reg [31:0] REG_427; // @[Hold.scala 89:18]
  reg [31:0] REG_428; // @[Hold.scala 89:18]
  reg [31:0] REG_429; // @[Hold.scala 89:18]
  reg [31:0] REG_430; // @[Hold.scala 89:18]
  reg [31:0] REG_431; // @[Hold.scala 89:18]
  reg [31:0] REG_432; // @[Hold.scala 89:18]
  reg [31:0] REG_433; // @[Hold.scala 89:18]
  reg [31:0] REG_434; // @[Hold.scala 89:18]
  reg [31:0] REG_435; // @[Hold.scala 89:18]
  reg [31:0] REG_436; // @[Hold.scala 89:18]
  reg [31:0] REG_437; // @[Hold.scala 89:18]
  reg [31:0] REG_438; // @[Hold.scala 89:18]
  reg [31:0] REG_439; // @[Hold.scala 89:18]
  reg [31:0] REG_440; // @[Hold.scala 89:18]
  reg [31:0] REG_441; // @[Hold.scala 89:18]
  reg [31:0] REG_442; // @[Hold.scala 89:18]
  reg [31:0] REG_443; // @[Hold.scala 89:18]
  reg [31:0] REG_444; // @[Hold.scala 89:18]
  reg [31:0] REG_445; // @[Hold.scala 89:18]
  reg [31:0] REG_446; // @[Hold.scala 89:18]
  reg [31:0] REG_447; // @[Hold.scala 89:18]
  reg [31:0] REG_448; // @[Hold.scala 89:18]
  reg [31:0] REG_449; // @[Hold.scala 89:18]
  reg [31:0] REG_450; // @[Hold.scala 89:18]
  reg [31:0] REG_451; // @[Hold.scala 89:18]
  reg [31:0] REG_452; // @[Hold.scala 89:18]
  reg [31:0] REG_453; // @[Hold.scala 89:18]
  reg [31:0] REG_454; // @[Hold.scala 89:18]
  reg [31:0] REG_455; // @[Hold.scala 89:18]
  reg [31:0] REG_456; // @[Hold.scala 89:18]
  reg [31:0] REG_457; // @[Hold.scala 89:18]
  reg [31:0] REG_458; // @[Hold.scala 89:18]
  reg [31:0] REG_459; // @[Hold.scala 89:18]
  reg [31:0] REG_460; // @[Hold.scala 89:18]
  reg [31:0] REG_461; // @[Hold.scala 89:18]
  reg [31:0] REG_462; // @[Hold.scala 89:18]
  reg [31:0] REG_463; // @[Hold.scala 89:18]
  reg [31:0] REG_464; // @[Hold.scala 89:18]
  reg [31:0] REG_465; // @[Hold.scala 89:18]
  reg [31:0] REG_466; // @[Hold.scala 89:18]
  reg [31:0] REG_467; // @[Hold.scala 89:18]
  reg [31:0] REG_468; // @[Hold.scala 89:18]
  reg [31:0] REG_469; // @[Hold.scala 89:18]
  reg [31:0] REG_470; // @[Hold.scala 89:18]
  reg [31:0] REG_471; // @[Hold.scala 89:18]
  reg [31:0] REG_472; // @[Hold.scala 89:18]
  reg [31:0] REG_473; // @[Hold.scala 89:18]
  reg [31:0] REG_474; // @[Hold.scala 89:18]
  reg [31:0] REG_475; // @[Hold.scala 89:18]
  reg [31:0] REG_476; // @[Hold.scala 89:18]
  reg [31:0] REG_477; // @[Hold.scala 89:18]
  reg [31:0] REG_478; // @[Hold.scala 89:18]
  reg [31:0] REG_479; // @[Hold.scala 89:18]
  reg [31:0] REG_480; // @[Hold.scala 89:18]
  reg [31:0] REG_481; // @[Hold.scala 89:18]
  reg [31:0] REG_482; // @[Hold.scala 89:18]
  reg [31:0] REG_483; // @[Hold.scala 89:18]
  reg [31:0] REG_484; // @[Hold.scala 89:18]
  reg [31:0] REG_485; // @[Hold.scala 89:18]
  reg [31:0] REG_486; // @[Hold.scala 89:18]
  reg [31:0] REG_487; // @[Hold.scala 89:18]
  reg [31:0] REG_488; // @[Hold.scala 89:18]
  reg [31:0] REG_489; // @[Hold.scala 89:18]
  reg [31:0] REG_490; // @[Hold.scala 89:18]
  reg [31:0] REG_491; // @[Hold.scala 89:18]
  reg [31:0] REG_492; // @[Hold.scala 89:18]
  reg [31:0] REG_493; // @[Hold.scala 89:18]
  reg [31:0] REG_494; // @[Hold.scala 89:18]
  reg [31:0] REG_495; // @[Hold.scala 89:18]
  reg [31:0] REG_496; // @[Hold.scala 89:18]
  reg [31:0] REG_497; // @[Hold.scala 89:18]
  reg [31:0] REG_498; // @[Hold.scala 89:18]
  reg [31:0] REG_499; // @[Hold.scala 89:18]
  reg [31:0] REG_500; // @[Hold.scala 89:18]
  reg [31:0] REG_501; // @[Hold.scala 89:18]
  reg [31:0] REG_502; // @[Hold.scala 89:18]
  reg [31:0] REG_503; // @[Hold.scala 89:18]
  reg [31:0] REG_504; // @[Hold.scala 89:18]
  reg [31:0] REG_505; // @[Hold.scala 89:18]
  reg [31:0] REG_506; // @[Hold.scala 89:18]
  reg [31:0] REG_507; // @[Hold.scala 89:18]
  reg [31:0] REG_508; // @[Hold.scala 89:18]
  reg [31:0] REG_509; // @[Hold.scala 89:18]
  reg [31:0] REG_510; // @[Hold.scala 89:18]
  reg [31:0] REG_511; // @[Hold.scala 89:18]
  reg [31:0] REG_512; // @[Hold.scala 89:18]
  reg [31:0] REG_513; // @[Hold.scala 89:18]
  reg [31:0] REG_514; // @[Hold.scala 89:18]
  reg [31:0] REG_515; // @[Hold.scala 89:18]
  reg [31:0] REG_516; // @[Hold.scala 89:18]
  reg [31:0] REG_517; // @[Hold.scala 89:18]
  reg [31:0] REG_518; // @[Hold.scala 89:18]
  reg [31:0] REG_519; // @[Hold.scala 89:18]
  reg [31:0] REG_520; // @[Hold.scala 89:18]
  reg [31:0] REG_521; // @[Hold.scala 89:18]
  reg [31:0] REG_522; // @[Hold.scala 89:18]
  reg [31:0] REG_523; // @[Hold.scala 89:18]
  reg [31:0] REG_524; // @[Hold.scala 89:18]
  reg [31:0] REG_525; // @[Hold.scala 89:18]
  reg [31:0] REG_526; // @[Hold.scala 89:18]
  reg [31:0] REG_527; // @[Hold.scala 89:18]
  reg [31:0] REG_528; // @[Hold.scala 89:18]
  reg [31:0] REG_529; // @[Hold.scala 89:18]
  reg [31:0] REG_530; // @[Hold.scala 89:18]
  reg [31:0] REG_531; // @[Hold.scala 89:18]
  reg [31:0] REG_532; // @[Hold.scala 89:18]
  reg [31:0] REG_533; // @[Hold.scala 89:18]
  reg [31:0] REG_534; // @[Hold.scala 89:18]
  reg [31:0] REG_535; // @[Hold.scala 89:18]
  reg [31:0] REG_536; // @[Hold.scala 89:18]
  reg [31:0] REG_537; // @[Hold.scala 89:18]
  reg [31:0] REG_538; // @[Hold.scala 89:18]
  reg [31:0] REG_539; // @[Hold.scala 89:18]
  reg [31:0] REG_540; // @[Hold.scala 89:18]
  reg [31:0] REG_541; // @[Hold.scala 89:18]
  reg [31:0] REG_542; // @[Hold.scala 89:18]
  reg [31:0] REG_543; // @[Hold.scala 89:18]
  reg [31:0] REG_544; // @[Hold.scala 89:18]
  reg [31:0] REG_545; // @[Hold.scala 89:18]
  reg [31:0] REG_546; // @[Hold.scala 89:18]
  reg [31:0] REG_547; // @[Hold.scala 89:18]
  reg [31:0] REG_548; // @[Hold.scala 89:18]
  reg [31:0] REG_549; // @[Hold.scala 89:18]
  reg [31:0] REG_550; // @[Hold.scala 89:18]
  reg [31:0] REG_551; // @[Hold.scala 89:18]
  reg [31:0] REG_552; // @[Hold.scala 89:18]
  reg [31:0] REG_553; // @[Hold.scala 89:18]
  reg [31:0] REG_554; // @[Hold.scala 89:18]
  reg [31:0] REG_555; // @[Hold.scala 89:18]
  reg [31:0] REG_556; // @[Hold.scala 89:18]
  reg [31:0] REG_557; // @[Hold.scala 89:18]
  reg [31:0] REG_558; // @[Hold.scala 89:18]
  reg [31:0] REG_559; // @[Hold.scala 89:18]
  reg [31:0] REG_560; // @[Hold.scala 89:18]
  reg [31:0] REG_561; // @[Hold.scala 89:18]
  reg [31:0] REG_562; // @[Hold.scala 89:18]
  reg [31:0] REG_563; // @[Hold.scala 89:18]
  reg [31:0] REG_564; // @[Hold.scala 89:18]
  reg [31:0] REG_565; // @[Hold.scala 89:18]
  reg [31:0] REG_566; // @[Hold.scala 89:18]
  reg [31:0] REG_567; // @[Hold.scala 89:18]
  reg [31:0] REG_568; // @[Hold.scala 89:18]
  reg [31:0] REG_569; // @[Hold.scala 89:18]
  reg [31:0] REG_570; // @[Hold.scala 89:18]
  reg [31:0] REG_571; // @[Hold.scala 89:18]
  reg [31:0] REG_572; // @[Hold.scala 89:18]
  reg [31:0] REG_573; // @[Hold.scala 89:18]
  reg [31:0] REG_574; // @[Hold.scala 89:18]
  reg [31:0] REG_575; // @[Hold.scala 89:18]
  reg [31:0] REG_576; // @[Hold.scala 89:18]
  reg [31:0] REG_577; // @[Hold.scala 89:18]
  reg [31:0] REG_578; // @[Hold.scala 89:18]
  reg [31:0] REG_579; // @[Hold.scala 89:18]
  reg [31:0] REG_580; // @[Hold.scala 89:18]
  reg [31:0] REG_581; // @[Hold.scala 89:18]
  reg [31:0] REG_582; // @[Hold.scala 89:18]
  reg [31:0] REG_583; // @[Hold.scala 89:18]
  reg [31:0] REG_584; // @[Hold.scala 89:18]
  reg [31:0] REG_585; // @[Hold.scala 89:18]
  reg [31:0] REG_586; // @[Hold.scala 89:18]
  reg [31:0] REG_587; // @[Hold.scala 89:18]
  reg [31:0] REG_588; // @[Hold.scala 89:18]
  reg [31:0] REG_589; // @[Hold.scala 89:18]
  reg [31:0] REG_590; // @[Hold.scala 89:18]
  reg [31:0] REG_591; // @[Hold.scala 89:18]
  reg [31:0] REG_592; // @[Hold.scala 89:18]
  reg [31:0] REG_593; // @[Hold.scala 89:18]
  reg [31:0] REG_594; // @[Hold.scala 89:18]
  reg [31:0] REG_595; // @[Hold.scala 89:18]
  reg [31:0] REG_596; // @[Hold.scala 89:18]
  reg [31:0] REG_597; // @[Hold.scala 89:18]
  reg [31:0] REG_598; // @[Hold.scala 89:18]
  reg [31:0] REG_599; // @[Hold.scala 89:18]
  reg [31:0] REG_600; // @[Hold.scala 89:18]
  reg [31:0] REG_601; // @[Hold.scala 89:18]
  reg [31:0] REG_602; // @[Hold.scala 89:18]
  reg [31:0] REG_603; // @[Hold.scala 89:18]
  reg [31:0] REG_604; // @[Hold.scala 89:18]
  reg [31:0] REG_605; // @[Hold.scala 89:18]
  reg [31:0] REG_606; // @[Hold.scala 89:18]
  reg [31:0] REG_607; // @[Hold.scala 89:18]
  reg [31:0] REG_608; // @[Hold.scala 89:18]
  reg [31:0] REG_609; // @[Hold.scala 89:18]
  reg [31:0] REG_610; // @[Hold.scala 89:18]
  reg [31:0] REG_611; // @[Hold.scala 89:18]
  reg [31:0] REG_612; // @[Hold.scala 89:18]
  reg [31:0] REG_613; // @[Hold.scala 89:18]
  reg [31:0] REG_614; // @[Hold.scala 89:18]
  reg [31:0] REG_615; // @[Hold.scala 89:18]
  reg [31:0] REG_616; // @[Hold.scala 89:18]
  reg [31:0] REG_617; // @[Hold.scala 89:18]
  reg [31:0] REG_618; // @[Hold.scala 89:18]
  reg [31:0] REG_619; // @[Hold.scala 89:18]
  reg [31:0] REG_620; // @[Hold.scala 89:18]
  reg [31:0] REG_621; // @[Hold.scala 89:18]
  reg [31:0] REG_622; // @[Hold.scala 89:18]
  reg [31:0] REG_623; // @[Hold.scala 89:18]
  reg [31:0] REG_624; // @[Hold.scala 89:18]
  reg [31:0] REG_625; // @[Hold.scala 89:18]
  reg [31:0] REG_626; // @[Hold.scala 89:18]
  reg [31:0] REG_627; // @[Hold.scala 89:18]
  reg [31:0] REG_628; // @[Hold.scala 89:18]
  reg [31:0] REG_629; // @[Hold.scala 89:18]
  reg [31:0] REG_630; // @[Hold.scala 89:18]
  reg [31:0] REG_631; // @[Hold.scala 89:18]
  reg [31:0] REG_632; // @[Hold.scala 89:18]
  reg [31:0] REG_633; // @[Hold.scala 89:18]
  reg [31:0] REG_634; // @[Hold.scala 89:18]
  reg [31:0] REG_635; // @[Hold.scala 89:18]
  reg [31:0] REG_636; // @[Hold.scala 89:18]
  reg [31:0] REG_637; // @[Hold.scala 89:18]
  reg [31:0] REG_638; // @[Hold.scala 89:18]
  reg [31:0] REG_639; // @[Hold.scala 89:18]
  reg [31:0] REG_640; // @[Hold.scala 89:18]
  reg [31:0] REG_641; // @[Hold.scala 89:18]
  reg [31:0] REG_642; // @[Hold.scala 89:18]
  reg [31:0] REG_643; // @[Hold.scala 89:18]
  reg [31:0] REG_644; // @[Hold.scala 89:18]
  reg [31:0] REG_645; // @[Hold.scala 89:18]
  reg [31:0] REG_646; // @[Hold.scala 89:18]
  reg [31:0] REG_647; // @[Hold.scala 89:18]
  reg [31:0] REG_648; // @[Hold.scala 89:18]
  reg [31:0] REG_649; // @[Hold.scala 89:18]
  reg [31:0] REG_650; // @[Hold.scala 89:18]
  reg [31:0] REG_651; // @[Hold.scala 89:18]
  reg [31:0] REG_652; // @[Hold.scala 89:18]
  reg [31:0] REG_653; // @[Hold.scala 89:18]
  reg [31:0] REG_654; // @[Hold.scala 89:18]
  reg [31:0] REG_655; // @[Hold.scala 89:18]
  reg [31:0] REG_656; // @[Hold.scala 89:18]
  reg [31:0] REG_657; // @[Hold.scala 89:18]
  reg [31:0] REG_658; // @[Hold.scala 89:18]
  reg [31:0] REG_659; // @[Hold.scala 89:18]
  reg [31:0] REG_660; // @[Hold.scala 89:18]
  reg [31:0] REG_661; // @[Hold.scala 89:18]
  reg [31:0] REG_662; // @[Hold.scala 89:18]
  reg [31:0] REG_663; // @[Hold.scala 89:18]
  reg [31:0] REG_664; // @[Hold.scala 89:18]
  reg [31:0] REG_665; // @[Hold.scala 89:18]
  reg [31:0] REG_666; // @[Hold.scala 89:18]
  reg [31:0] REG_667; // @[Hold.scala 89:18]
  reg [31:0] REG_668; // @[Hold.scala 89:18]
  reg [31:0] REG_669; // @[Hold.scala 89:18]
  reg [31:0] REG_670; // @[Hold.scala 89:18]
  reg [31:0] REG_671; // @[Hold.scala 89:18]
  reg [31:0] REG_672; // @[Hold.scala 89:18]
  reg [31:0] REG_673; // @[Hold.scala 89:18]
  reg [31:0] REG_674; // @[Hold.scala 89:18]
  reg [31:0] REG_675; // @[Hold.scala 89:18]
  reg [31:0] REG_676; // @[Hold.scala 89:18]
  reg [31:0] REG_677; // @[Hold.scala 89:18]
  reg [31:0] REG_678; // @[Hold.scala 89:18]
  reg [31:0] REG_679; // @[Hold.scala 89:18]
  reg [31:0] REG_680; // @[Hold.scala 89:18]
  reg [31:0] REG_681; // @[Hold.scala 89:18]
  reg [31:0] REG_682; // @[Hold.scala 89:18]
  reg [31:0] REG_683; // @[Hold.scala 89:18]
  reg [31:0] REG_684; // @[Hold.scala 89:18]
  reg [31:0] REG_685; // @[Hold.scala 89:18]
  reg [31:0] REG_686; // @[Hold.scala 89:18]
  reg [31:0] REG_687; // @[Hold.scala 89:18]
  reg [31:0] REG_688; // @[Hold.scala 89:18]
  reg [31:0] REG_689; // @[Hold.scala 89:18]
  reg [31:0] REG_690; // @[Hold.scala 89:18]
  reg [31:0] REG_691; // @[Hold.scala 89:18]
  reg [31:0] REG_692; // @[Hold.scala 89:18]
  reg [31:0] REG_693; // @[Hold.scala 89:18]
  reg [31:0] REG_694; // @[Hold.scala 89:18]
  reg [31:0] REG_695; // @[Hold.scala 89:18]
  reg [31:0] REG_696; // @[Hold.scala 89:18]
  reg [31:0] REG_697; // @[Hold.scala 89:18]
  reg [31:0] REG_698; // @[Hold.scala 89:18]
  reg [31:0] REG_699; // @[Hold.scala 89:18]
  reg [31:0] REG_700; // @[Hold.scala 89:18]
  reg [31:0] REG_701; // @[Hold.scala 89:18]
  reg [31:0] REG_702; // @[Hold.scala 89:18]
  reg [31:0] REG_703; // @[Hold.scala 89:18]
  reg [31:0] REG_704; // @[Hold.scala 89:18]
  reg [31:0] REG_705; // @[Hold.scala 89:18]
  reg [31:0] REG_706; // @[Hold.scala 89:18]
  reg [31:0] REG_707; // @[Hold.scala 89:18]
  reg [31:0] REG_708; // @[Hold.scala 89:18]
  reg [31:0] REG_709; // @[Hold.scala 89:18]
  reg [31:0] REG_710; // @[Hold.scala 89:18]
  reg [31:0] REG_711; // @[Hold.scala 89:18]
  reg [31:0] REG_712; // @[Hold.scala 89:18]
  reg [31:0] REG_713; // @[Hold.scala 89:18]
  reg [31:0] REG_714; // @[Hold.scala 89:18]
  reg [31:0] REG_715; // @[Hold.scala 89:18]
  reg [31:0] REG_716; // @[Hold.scala 89:18]
  reg [31:0] REG_717; // @[Hold.scala 89:18]
  reg [31:0] REG_718; // @[Hold.scala 89:18]
  reg [31:0] REG_719; // @[Hold.scala 89:18]
  reg [31:0] REG_720; // @[Hold.scala 89:18]
  reg [31:0] REG_721; // @[Hold.scala 89:18]
  reg [31:0] REG_722; // @[Hold.scala 89:18]
  reg [31:0] REG_723; // @[Hold.scala 89:18]
  reg [31:0] REG_724; // @[Hold.scala 89:18]
  reg [31:0] REG_725; // @[Hold.scala 89:18]
  reg [31:0] REG_726; // @[Hold.scala 89:18]
  reg [31:0] REG_727; // @[Hold.scala 89:18]
  reg [31:0] REG_728; // @[Hold.scala 89:18]
  reg [31:0] REG_729; // @[Hold.scala 89:18]
  reg [31:0] REG_730; // @[Hold.scala 89:18]
  reg [31:0] REG_731; // @[Hold.scala 89:18]
  reg [31:0] REG_732; // @[Hold.scala 89:18]
  reg [31:0] REG_733; // @[Hold.scala 89:18]
  reg [31:0] REG_734; // @[Hold.scala 89:18]
  reg [31:0] REG_735; // @[Hold.scala 89:18]
  reg [31:0] REG_736; // @[Hold.scala 89:18]
  reg [31:0] REG_737; // @[Hold.scala 89:18]
  reg [31:0] REG_738; // @[Hold.scala 89:18]
  reg [31:0] REG_739; // @[Hold.scala 89:18]
  reg [31:0] REG_740; // @[Hold.scala 89:18]
  reg [31:0] REG_741; // @[Hold.scala 89:18]
  reg [31:0] REG_742; // @[Hold.scala 89:18]
  reg [31:0] REG_743; // @[Hold.scala 89:18]
  reg [31:0] REG_744; // @[Hold.scala 89:18]
  reg [31:0] REG_745; // @[Hold.scala 89:18]
  reg [31:0] REG_746; // @[Hold.scala 89:18]
  reg [31:0] REG_747; // @[Hold.scala 89:18]
  reg [31:0] REG_748; // @[Hold.scala 89:18]
  reg [31:0] REG_749; // @[Hold.scala 89:18]
  reg [31:0] REG_750; // @[Hold.scala 89:18]
  reg [31:0] REG_751; // @[Hold.scala 89:18]
  reg [31:0] REG_752; // @[Hold.scala 89:18]
  reg [31:0] REG_753; // @[Hold.scala 89:18]
  reg [31:0] REG_754; // @[Hold.scala 89:18]
  reg [31:0] REG_755; // @[Hold.scala 89:18]
  reg [31:0] REG_756; // @[Hold.scala 89:18]
  reg [31:0] REG_757; // @[Hold.scala 89:18]
  reg [31:0] REG_758; // @[Hold.scala 89:18]
  reg [31:0] REG_759; // @[Hold.scala 89:18]
  reg [31:0] REG_760; // @[Hold.scala 89:18]
  reg [31:0] REG_761; // @[Hold.scala 89:18]
  reg [31:0] REG_762; // @[Hold.scala 89:18]
  reg [31:0] REG_763; // @[Hold.scala 89:18]
  reg [31:0] REG_764; // @[Hold.scala 89:18]
  reg [31:0] REG_765; // @[Hold.scala 89:18]
  reg [31:0] REG_766; // @[Hold.scala 89:18]
  reg [31:0] REG_767; // @[Hold.scala 89:18]
  reg [31:0] REG_768; // @[Hold.scala 89:18]
  reg [31:0] REG_769; // @[Hold.scala 89:18]
  reg [31:0] REG_770; // @[Hold.scala 89:18]
  reg [31:0] REG_771; // @[Hold.scala 89:18]
  reg [31:0] REG_772; // @[Hold.scala 89:18]
  reg [31:0] REG_773; // @[Hold.scala 89:18]
  reg [31:0] REG_774; // @[Hold.scala 89:18]
  reg [31:0] REG_775; // @[Hold.scala 89:18]
  reg [31:0] REG_776; // @[Hold.scala 89:18]
  reg [31:0] REG_777; // @[Hold.scala 89:18]
  reg [31:0] REG_778; // @[Hold.scala 89:18]
  reg [31:0] REG_779; // @[Hold.scala 89:18]
  reg [31:0] REG_780; // @[Hold.scala 89:18]
  reg [31:0] REG_781; // @[Hold.scala 89:18]
  reg [31:0] REG_782; // @[Hold.scala 89:18]
  reg [31:0] REG_783; // @[Hold.scala 89:18]
  reg [31:0] REG_784; // @[Hold.scala 89:18]
  reg [31:0] REG_785; // @[Hold.scala 89:18]
  reg [31:0] REG_786; // @[Hold.scala 89:18]
  reg [31:0] REG_787; // @[Hold.scala 89:18]
  reg [31:0] REG_788; // @[Hold.scala 89:18]
  reg [31:0] REG_789; // @[Hold.scala 89:18]
  reg [31:0] REG_790; // @[Hold.scala 89:18]
  reg [31:0] REG_791; // @[Hold.scala 89:18]
  reg [31:0] REG_792; // @[Hold.scala 89:18]
  reg [31:0] REG_793; // @[Hold.scala 89:18]
  reg [31:0] REG_794; // @[Hold.scala 89:18]
  reg [31:0] REG_795; // @[Hold.scala 89:18]
  reg [31:0] REG_796; // @[Hold.scala 89:18]
  reg [31:0] REG_797; // @[Hold.scala 89:18]
  reg [31:0] REG_798; // @[Hold.scala 89:18]
  reg [31:0] REG_799; // @[Hold.scala 89:18]
  reg [31:0] REG_800; // @[Hold.scala 89:18]
  reg [31:0] REG_801; // @[Hold.scala 89:18]
  reg [31:0] REG_802; // @[Hold.scala 89:18]
  reg [31:0] REG_803; // @[Hold.scala 89:18]
  reg [31:0] REG_804; // @[Hold.scala 89:18]
  reg [31:0] REG_805; // @[Hold.scala 89:18]
  reg [31:0] REG_806; // @[Hold.scala 89:18]
  reg [31:0] REG_807; // @[Hold.scala 89:18]
  reg [31:0] REG_808; // @[Hold.scala 89:18]
  reg [31:0] REG_809; // @[Hold.scala 89:18]
  reg [31:0] REG_810; // @[Hold.scala 89:18]
  reg [31:0] REG_811; // @[Hold.scala 89:18]
  reg [31:0] REG_812; // @[Hold.scala 89:18]
  reg [31:0] REG_813; // @[Hold.scala 89:18]
  reg [31:0] REG_814; // @[Hold.scala 89:18]
  reg [31:0] REG_815; // @[Hold.scala 89:18]
  reg [31:0] REG_816; // @[Hold.scala 89:18]
  reg [31:0] REG_817; // @[Hold.scala 89:18]
  reg [31:0] REG_818; // @[Hold.scala 89:18]
  reg [31:0] REG_819; // @[Hold.scala 89:18]
  reg [31:0] REG_820; // @[Hold.scala 89:18]
  reg [31:0] REG_821; // @[Hold.scala 89:18]
  reg [31:0] REG_822; // @[Hold.scala 89:18]
  reg [31:0] REG_823; // @[Hold.scala 89:18]
  reg [31:0] REG_824; // @[Hold.scala 89:18]
  reg [31:0] REG_825; // @[Hold.scala 89:18]
  reg [31:0] REG_826; // @[Hold.scala 89:18]
  reg [31:0] REG_827; // @[Hold.scala 89:18]
  reg [31:0] REG_828; // @[Hold.scala 89:18]
  reg [31:0] REG_829; // @[Hold.scala 89:18]
  reg [31:0] REG_830; // @[Hold.scala 89:18]
  reg [31:0] REG_831; // @[Hold.scala 89:18]
  reg [31:0] REG_832; // @[Hold.scala 89:18]
  reg [31:0] REG_833; // @[Hold.scala 89:18]
  reg [31:0] REG_834; // @[Hold.scala 89:18]
  reg [31:0] REG_835; // @[Hold.scala 89:18]
  reg [31:0] REG_836; // @[Hold.scala 89:18]
  reg [31:0] REG_837; // @[Hold.scala 89:18]
  reg [31:0] REG_838; // @[Hold.scala 89:18]
  reg [31:0] REG_839; // @[Hold.scala 89:18]
  reg [31:0] REG_840; // @[Hold.scala 89:18]
  reg [31:0] REG_841; // @[Hold.scala 89:18]
  reg [31:0] REG_842; // @[Hold.scala 89:18]
  reg [31:0] REG_843; // @[Hold.scala 89:18]
  reg [31:0] REG_844; // @[Hold.scala 89:18]
  reg [31:0] REG_845; // @[Hold.scala 89:18]
  reg [31:0] REG_846; // @[Hold.scala 89:18]
  reg [31:0] REG_847; // @[Hold.scala 89:18]
  reg [31:0] REG_848; // @[Hold.scala 89:18]
  reg [31:0] REG_849; // @[Hold.scala 89:18]
  reg [31:0] REG_850; // @[Hold.scala 89:18]
  reg [31:0] REG_851; // @[Hold.scala 89:18]
  reg [31:0] REG_852; // @[Hold.scala 89:18]
  reg [31:0] REG_853; // @[Hold.scala 89:18]
  reg [31:0] REG_854; // @[Hold.scala 89:18]
  reg [31:0] REG_855; // @[Hold.scala 89:18]
  reg [31:0] REG_856; // @[Hold.scala 89:18]
  reg [31:0] REG_857; // @[Hold.scala 89:18]
  reg [31:0] REG_858; // @[Hold.scala 89:18]
  reg [31:0] REG_859; // @[Hold.scala 89:18]
  reg [31:0] REG_860; // @[Hold.scala 89:18]
  reg [31:0] REG_861; // @[Hold.scala 89:18]
  reg [31:0] REG_862; // @[Hold.scala 89:18]
  reg [31:0] REG_863; // @[Hold.scala 89:18]
  reg [31:0] REG_864; // @[Hold.scala 89:18]
  reg [31:0] REG_865; // @[Hold.scala 89:18]
  reg [31:0] REG_866; // @[Hold.scala 89:18]
  reg [31:0] REG_867; // @[Hold.scala 89:18]
  reg [31:0] REG_868; // @[Hold.scala 89:18]
  reg [31:0] REG_869; // @[Hold.scala 89:18]
  reg [31:0] REG_870; // @[Hold.scala 89:18]
  reg [31:0] REG_871; // @[Hold.scala 89:18]
  reg [31:0] REG_872; // @[Hold.scala 89:18]
  reg [31:0] REG_873; // @[Hold.scala 89:18]
  reg [31:0] REG_874; // @[Hold.scala 89:18]
  reg [31:0] REG_875; // @[Hold.scala 89:18]
  reg [31:0] REG_876; // @[Hold.scala 89:18]
  reg [31:0] REG_877; // @[Hold.scala 89:18]
  reg [31:0] REG_878; // @[Hold.scala 89:18]
  reg [31:0] REG_879; // @[Hold.scala 89:18]
  reg [31:0] REG_880; // @[Hold.scala 89:18]
  reg [31:0] REG_881; // @[Hold.scala 89:18]
  reg [31:0] REG_882; // @[Hold.scala 89:18]
  reg [31:0] REG_883; // @[Hold.scala 89:18]
  reg [31:0] REG_884; // @[Hold.scala 89:18]
  reg [31:0] REG_885; // @[Hold.scala 89:18]
  reg [31:0] REG_886; // @[Hold.scala 89:18]
  reg [31:0] REG_887; // @[Hold.scala 89:18]
  reg [31:0] REG_888; // @[Hold.scala 89:18]
  reg [31:0] REG_889; // @[Hold.scala 89:18]
  reg [31:0] REG_890; // @[Hold.scala 89:18]
  reg [31:0] REG_891; // @[Hold.scala 89:18]
  reg [31:0] REG_892; // @[Hold.scala 89:18]
  reg [31:0] REG_893; // @[Hold.scala 89:18]
  reg [31:0] REG_894; // @[Hold.scala 89:18]
  reg [31:0] REG_895; // @[Hold.scala 89:18]
  reg [31:0] REG_896; // @[Hold.scala 89:18]
  reg [31:0] REG_897; // @[Hold.scala 89:18]
  reg [31:0] REG_898; // @[Hold.scala 89:18]
  reg [31:0] REG_899; // @[Hold.scala 89:18]
  reg [31:0] REG_900; // @[Hold.scala 89:18]
  reg [31:0] REG_901; // @[Hold.scala 89:18]
  reg [31:0] REG_902; // @[Hold.scala 89:18]
  reg [31:0] REG_903; // @[Hold.scala 89:18]
  reg [31:0] REG_904; // @[Hold.scala 89:18]
  reg [31:0] REG_905; // @[Hold.scala 89:18]
  reg [31:0] REG_906; // @[Hold.scala 89:18]
  reg [31:0] REG_907; // @[Hold.scala 89:18]
  reg [31:0] REG_908; // @[Hold.scala 89:18]
  reg [31:0] REG_909; // @[Hold.scala 89:18]
  reg [31:0] REG_910; // @[Hold.scala 89:18]
  reg [31:0] REG_911; // @[Hold.scala 89:18]
  reg [31:0] REG_912; // @[Hold.scala 89:18]
  reg [31:0] REG_913; // @[Hold.scala 89:18]
  reg [31:0] REG_914; // @[Hold.scala 89:18]
  reg [31:0] REG_915; // @[Hold.scala 89:18]
  reg [31:0] REG_916; // @[Hold.scala 89:18]
  reg [31:0] REG_917; // @[Hold.scala 89:18]
  reg [31:0] REG_918; // @[Hold.scala 89:18]
  reg [31:0] REG_919; // @[Hold.scala 89:18]
  reg [31:0] REG_920; // @[Hold.scala 89:18]
  reg [31:0] REG_921; // @[Hold.scala 89:18]
  reg [31:0] REG_922; // @[Hold.scala 89:18]
  reg [31:0] REG_923; // @[Hold.scala 89:18]
  reg [31:0] REG_924; // @[Hold.scala 89:18]
  reg [31:0] REG_925; // @[Hold.scala 89:18]
  reg [31:0] REG_926; // @[Hold.scala 89:18]
  reg [31:0] REG_927; // @[Hold.scala 89:18]
  reg [31:0] REG_928; // @[Hold.scala 89:18]
  reg [31:0] REG_929; // @[Hold.scala 89:18]
  reg [31:0] REG_930; // @[Hold.scala 89:18]
  reg [31:0] REG_931; // @[Hold.scala 89:18]
  reg [31:0] REG_932; // @[Hold.scala 89:18]
  reg [31:0] REG_933; // @[Hold.scala 89:18]
  reg [31:0] REG_934; // @[Hold.scala 89:18]
  reg [31:0] REG_935; // @[Hold.scala 89:18]
  reg [31:0] REG_936; // @[Hold.scala 89:18]
  reg [31:0] REG_937; // @[Hold.scala 89:18]
  reg [31:0] REG_938; // @[Hold.scala 89:18]
  reg [31:0] REG_939; // @[Hold.scala 89:18]
  reg [31:0] REG_940; // @[Hold.scala 89:18]
  reg [31:0] REG_941; // @[Hold.scala 89:18]
  reg [31:0] REG_942; // @[Hold.scala 89:18]
  reg [31:0] REG_943; // @[Hold.scala 89:18]
  reg [31:0] REG_944; // @[Hold.scala 89:18]
  reg [31:0] REG_945; // @[Hold.scala 89:18]
  reg [31:0] REG_946; // @[Hold.scala 89:18]
  reg [31:0] REG_947; // @[Hold.scala 89:18]
  reg [31:0] REG_948; // @[Hold.scala 89:18]
  reg [31:0] REG_949; // @[Hold.scala 89:18]
  reg [31:0] REG_950; // @[Hold.scala 89:18]
  reg [31:0] REG_951; // @[Hold.scala 89:18]
  reg [31:0] REG_952; // @[Hold.scala 89:18]
  reg [31:0] REG_953; // @[Hold.scala 89:18]
  reg [31:0] REG_954; // @[Hold.scala 89:18]
  reg [31:0] REG_955; // @[Hold.scala 89:18]
  reg [31:0] REG_956; // @[Hold.scala 89:18]
  reg [31:0] REG_957; // @[Hold.scala 89:18]
  reg [31:0] REG_958; // @[Hold.scala 89:18]
  reg [31:0] REG_959; // @[Hold.scala 89:18]
  reg [31:0] REG_960; // @[Hold.scala 89:18]
  reg [31:0] REG_961; // @[Hold.scala 89:18]
  reg [31:0] REG_962; // @[Hold.scala 89:18]
  reg [31:0] REG_963; // @[Hold.scala 89:18]
  reg [31:0] REG_964; // @[Hold.scala 89:18]
  reg [31:0] REG_965; // @[Hold.scala 89:18]
  reg [31:0] REG_966; // @[Hold.scala 89:18]
  reg [31:0] REG_967; // @[Hold.scala 89:18]
  reg [31:0] REG_968; // @[Hold.scala 89:18]
  reg [31:0] REG_969; // @[Hold.scala 89:18]
  reg [31:0] REG_970; // @[Hold.scala 89:18]
  reg [31:0] REG_971; // @[Hold.scala 89:18]
  reg [31:0] REG_972; // @[Hold.scala 89:18]
  reg [31:0] REG_973; // @[Hold.scala 89:18]
  reg [31:0] REG_974; // @[Hold.scala 89:18]
  reg [31:0] REG_975; // @[Hold.scala 89:18]
  reg [31:0] REG_976; // @[Hold.scala 89:18]
  reg [31:0] REG_977; // @[Hold.scala 89:18]
  reg [31:0] REG_978; // @[Hold.scala 89:18]
  reg [31:0] REG_979; // @[Hold.scala 89:18]
  reg [31:0] REG_980; // @[Hold.scala 89:18]
  reg [31:0] REG_981; // @[Hold.scala 89:18]
  reg [31:0] REG_982; // @[Hold.scala 89:18]
  reg [31:0] REG_983; // @[Hold.scala 89:18]
  reg [31:0] REG_984; // @[Hold.scala 89:18]
  reg [31:0] REG_985; // @[Hold.scala 89:18]
  reg [31:0] REG_986; // @[Hold.scala 89:18]
  reg [31:0] REG_987; // @[Hold.scala 89:18]
  reg [31:0] REG_988; // @[Hold.scala 89:18]
  reg [31:0] REG_989; // @[Hold.scala 89:18]
  reg [31:0] REG_990; // @[Hold.scala 89:18]
  reg [31:0] REG_991; // @[Hold.scala 89:18]
  reg [31:0] REG_992; // @[Hold.scala 89:18]
  reg [31:0] REG_993; // @[Hold.scala 89:18]
  reg [31:0] REG_994; // @[Hold.scala 89:18]
  reg [31:0] REG_995; // @[Hold.scala 89:18]
  reg [31:0] REG_996; // @[Hold.scala 89:18]
  reg [31:0] REG_997; // @[Hold.scala 89:18]
  reg [31:0] REG_998; // @[Hold.scala 89:18]
  reg [31:0] out; // @[Hold.scala 89:18]
  assign io_out = out; // @[Hold.scala 91:10]
  always @(posedge clock) begin
    REG <= io_in; // @[Hold.scala 89:18]
    REG_1 <= REG; // @[Hold.scala 89:18]
    REG_2 <= REG_1; // @[Hold.scala 89:18]
    REG_3 <= REG_2; // @[Hold.scala 89:18]
    REG_4 <= REG_3; // @[Hold.scala 89:18]
    REG_5 <= REG_4; // @[Hold.scala 89:18]
    REG_6 <= REG_5; // @[Hold.scala 89:18]
    REG_7 <= REG_6; // @[Hold.scala 89:18]
    REG_8 <= REG_7; // @[Hold.scala 89:18]
    REG_9 <= REG_8; // @[Hold.scala 89:18]
    REG_10 <= REG_9; // @[Hold.scala 89:18]
    REG_11 <= REG_10; // @[Hold.scala 89:18]
    REG_12 <= REG_11; // @[Hold.scala 89:18]
    REG_13 <= REG_12; // @[Hold.scala 89:18]
    REG_14 <= REG_13; // @[Hold.scala 89:18]
    REG_15 <= REG_14; // @[Hold.scala 89:18]
    REG_16 <= REG_15; // @[Hold.scala 89:18]
    REG_17 <= REG_16; // @[Hold.scala 89:18]
    REG_18 <= REG_17; // @[Hold.scala 89:18]
    REG_19 <= REG_18; // @[Hold.scala 89:18]
    REG_20 <= REG_19; // @[Hold.scala 89:18]
    REG_21 <= REG_20; // @[Hold.scala 89:18]
    REG_22 <= REG_21; // @[Hold.scala 89:18]
    REG_23 <= REG_22; // @[Hold.scala 89:18]
    REG_24 <= REG_23; // @[Hold.scala 89:18]
    REG_25 <= REG_24; // @[Hold.scala 89:18]
    REG_26 <= REG_25; // @[Hold.scala 89:18]
    REG_27 <= REG_26; // @[Hold.scala 89:18]
    REG_28 <= REG_27; // @[Hold.scala 89:18]
    REG_29 <= REG_28; // @[Hold.scala 89:18]
    REG_30 <= REG_29; // @[Hold.scala 89:18]
    REG_31 <= REG_30; // @[Hold.scala 89:18]
    REG_32 <= REG_31; // @[Hold.scala 89:18]
    REG_33 <= REG_32; // @[Hold.scala 89:18]
    REG_34 <= REG_33; // @[Hold.scala 89:18]
    REG_35 <= REG_34; // @[Hold.scala 89:18]
    REG_36 <= REG_35; // @[Hold.scala 89:18]
    REG_37 <= REG_36; // @[Hold.scala 89:18]
    REG_38 <= REG_37; // @[Hold.scala 89:18]
    REG_39 <= REG_38; // @[Hold.scala 89:18]
    REG_40 <= REG_39; // @[Hold.scala 89:18]
    REG_41 <= REG_40; // @[Hold.scala 89:18]
    REG_42 <= REG_41; // @[Hold.scala 89:18]
    REG_43 <= REG_42; // @[Hold.scala 89:18]
    REG_44 <= REG_43; // @[Hold.scala 89:18]
    REG_45 <= REG_44; // @[Hold.scala 89:18]
    REG_46 <= REG_45; // @[Hold.scala 89:18]
    REG_47 <= REG_46; // @[Hold.scala 89:18]
    REG_48 <= REG_47; // @[Hold.scala 89:18]
    REG_49 <= REG_48; // @[Hold.scala 89:18]
    REG_50 <= REG_49; // @[Hold.scala 89:18]
    REG_51 <= REG_50; // @[Hold.scala 89:18]
    REG_52 <= REG_51; // @[Hold.scala 89:18]
    REG_53 <= REG_52; // @[Hold.scala 89:18]
    REG_54 <= REG_53; // @[Hold.scala 89:18]
    REG_55 <= REG_54; // @[Hold.scala 89:18]
    REG_56 <= REG_55; // @[Hold.scala 89:18]
    REG_57 <= REG_56; // @[Hold.scala 89:18]
    REG_58 <= REG_57; // @[Hold.scala 89:18]
    REG_59 <= REG_58; // @[Hold.scala 89:18]
    REG_60 <= REG_59; // @[Hold.scala 89:18]
    REG_61 <= REG_60; // @[Hold.scala 89:18]
    REG_62 <= REG_61; // @[Hold.scala 89:18]
    REG_63 <= REG_62; // @[Hold.scala 89:18]
    REG_64 <= REG_63; // @[Hold.scala 89:18]
    REG_65 <= REG_64; // @[Hold.scala 89:18]
    REG_66 <= REG_65; // @[Hold.scala 89:18]
    REG_67 <= REG_66; // @[Hold.scala 89:18]
    REG_68 <= REG_67; // @[Hold.scala 89:18]
    REG_69 <= REG_68; // @[Hold.scala 89:18]
    REG_70 <= REG_69; // @[Hold.scala 89:18]
    REG_71 <= REG_70; // @[Hold.scala 89:18]
    REG_72 <= REG_71; // @[Hold.scala 89:18]
    REG_73 <= REG_72; // @[Hold.scala 89:18]
    REG_74 <= REG_73; // @[Hold.scala 89:18]
    REG_75 <= REG_74; // @[Hold.scala 89:18]
    REG_76 <= REG_75; // @[Hold.scala 89:18]
    REG_77 <= REG_76; // @[Hold.scala 89:18]
    REG_78 <= REG_77; // @[Hold.scala 89:18]
    REG_79 <= REG_78; // @[Hold.scala 89:18]
    REG_80 <= REG_79; // @[Hold.scala 89:18]
    REG_81 <= REG_80; // @[Hold.scala 89:18]
    REG_82 <= REG_81; // @[Hold.scala 89:18]
    REG_83 <= REG_82; // @[Hold.scala 89:18]
    REG_84 <= REG_83; // @[Hold.scala 89:18]
    REG_85 <= REG_84; // @[Hold.scala 89:18]
    REG_86 <= REG_85; // @[Hold.scala 89:18]
    REG_87 <= REG_86; // @[Hold.scala 89:18]
    REG_88 <= REG_87; // @[Hold.scala 89:18]
    REG_89 <= REG_88; // @[Hold.scala 89:18]
    REG_90 <= REG_89; // @[Hold.scala 89:18]
    REG_91 <= REG_90; // @[Hold.scala 89:18]
    REG_92 <= REG_91; // @[Hold.scala 89:18]
    REG_93 <= REG_92; // @[Hold.scala 89:18]
    REG_94 <= REG_93; // @[Hold.scala 89:18]
    REG_95 <= REG_94; // @[Hold.scala 89:18]
    REG_96 <= REG_95; // @[Hold.scala 89:18]
    REG_97 <= REG_96; // @[Hold.scala 89:18]
    REG_98 <= REG_97; // @[Hold.scala 89:18]
    REG_99 <= REG_98; // @[Hold.scala 89:18]
    REG_100 <= REG_99; // @[Hold.scala 89:18]
    REG_101 <= REG_100; // @[Hold.scala 89:18]
    REG_102 <= REG_101; // @[Hold.scala 89:18]
    REG_103 <= REG_102; // @[Hold.scala 89:18]
    REG_104 <= REG_103; // @[Hold.scala 89:18]
    REG_105 <= REG_104; // @[Hold.scala 89:18]
    REG_106 <= REG_105; // @[Hold.scala 89:18]
    REG_107 <= REG_106; // @[Hold.scala 89:18]
    REG_108 <= REG_107; // @[Hold.scala 89:18]
    REG_109 <= REG_108; // @[Hold.scala 89:18]
    REG_110 <= REG_109; // @[Hold.scala 89:18]
    REG_111 <= REG_110; // @[Hold.scala 89:18]
    REG_112 <= REG_111; // @[Hold.scala 89:18]
    REG_113 <= REG_112; // @[Hold.scala 89:18]
    REG_114 <= REG_113; // @[Hold.scala 89:18]
    REG_115 <= REG_114; // @[Hold.scala 89:18]
    REG_116 <= REG_115; // @[Hold.scala 89:18]
    REG_117 <= REG_116; // @[Hold.scala 89:18]
    REG_118 <= REG_117; // @[Hold.scala 89:18]
    REG_119 <= REG_118; // @[Hold.scala 89:18]
    REG_120 <= REG_119; // @[Hold.scala 89:18]
    REG_121 <= REG_120; // @[Hold.scala 89:18]
    REG_122 <= REG_121; // @[Hold.scala 89:18]
    REG_123 <= REG_122; // @[Hold.scala 89:18]
    REG_124 <= REG_123; // @[Hold.scala 89:18]
    REG_125 <= REG_124; // @[Hold.scala 89:18]
    REG_126 <= REG_125; // @[Hold.scala 89:18]
    REG_127 <= REG_126; // @[Hold.scala 89:18]
    REG_128 <= REG_127; // @[Hold.scala 89:18]
    REG_129 <= REG_128; // @[Hold.scala 89:18]
    REG_130 <= REG_129; // @[Hold.scala 89:18]
    REG_131 <= REG_130; // @[Hold.scala 89:18]
    REG_132 <= REG_131; // @[Hold.scala 89:18]
    REG_133 <= REG_132; // @[Hold.scala 89:18]
    REG_134 <= REG_133; // @[Hold.scala 89:18]
    REG_135 <= REG_134; // @[Hold.scala 89:18]
    REG_136 <= REG_135; // @[Hold.scala 89:18]
    REG_137 <= REG_136; // @[Hold.scala 89:18]
    REG_138 <= REG_137; // @[Hold.scala 89:18]
    REG_139 <= REG_138; // @[Hold.scala 89:18]
    REG_140 <= REG_139; // @[Hold.scala 89:18]
    REG_141 <= REG_140; // @[Hold.scala 89:18]
    REG_142 <= REG_141; // @[Hold.scala 89:18]
    REG_143 <= REG_142; // @[Hold.scala 89:18]
    REG_144 <= REG_143; // @[Hold.scala 89:18]
    REG_145 <= REG_144; // @[Hold.scala 89:18]
    REG_146 <= REG_145; // @[Hold.scala 89:18]
    REG_147 <= REG_146; // @[Hold.scala 89:18]
    REG_148 <= REG_147; // @[Hold.scala 89:18]
    REG_149 <= REG_148; // @[Hold.scala 89:18]
    REG_150 <= REG_149; // @[Hold.scala 89:18]
    REG_151 <= REG_150; // @[Hold.scala 89:18]
    REG_152 <= REG_151; // @[Hold.scala 89:18]
    REG_153 <= REG_152; // @[Hold.scala 89:18]
    REG_154 <= REG_153; // @[Hold.scala 89:18]
    REG_155 <= REG_154; // @[Hold.scala 89:18]
    REG_156 <= REG_155; // @[Hold.scala 89:18]
    REG_157 <= REG_156; // @[Hold.scala 89:18]
    REG_158 <= REG_157; // @[Hold.scala 89:18]
    REG_159 <= REG_158; // @[Hold.scala 89:18]
    REG_160 <= REG_159; // @[Hold.scala 89:18]
    REG_161 <= REG_160; // @[Hold.scala 89:18]
    REG_162 <= REG_161; // @[Hold.scala 89:18]
    REG_163 <= REG_162; // @[Hold.scala 89:18]
    REG_164 <= REG_163; // @[Hold.scala 89:18]
    REG_165 <= REG_164; // @[Hold.scala 89:18]
    REG_166 <= REG_165; // @[Hold.scala 89:18]
    REG_167 <= REG_166; // @[Hold.scala 89:18]
    REG_168 <= REG_167; // @[Hold.scala 89:18]
    REG_169 <= REG_168; // @[Hold.scala 89:18]
    REG_170 <= REG_169; // @[Hold.scala 89:18]
    REG_171 <= REG_170; // @[Hold.scala 89:18]
    REG_172 <= REG_171; // @[Hold.scala 89:18]
    REG_173 <= REG_172; // @[Hold.scala 89:18]
    REG_174 <= REG_173; // @[Hold.scala 89:18]
    REG_175 <= REG_174; // @[Hold.scala 89:18]
    REG_176 <= REG_175; // @[Hold.scala 89:18]
    REG_177 <= REG_176; // @[Hold.scala 89:18]
    REG_178 <= REG_177; // @[Hold.scala 89:18]
    REG_179 <= REG_178; // @[Hold.scala 89:18]
    REG_180 <= REG_179; // @[Hold.scala 89:18]
    REG_181 <= REG_180; // @[Hold.scala 89:18]
    REG_182 <= REG_181; // @[Hold.scala 89:18]
    REG_183 <= REG_182; // @[Hold.scala 89:18]
    REG_184 <= REG_183; // @[Hold.scala 89:18]
    REG_185 <= REG_184; // @[Hold.scala 89:18]
    REG_186 <= REG_185; // @[Hold.scala 89:18]
    REG_187 <= REG_186; // @[Hold.scala 89:18]
    REG_188 <= REG_187; // @[Hold.scala 89:18]
    REG_189 <= REG_188; // @[Hold.scala 89:18]
    REG_190 <= REG_189; // @[Hold.scala 89:18]
    REG_191 <= REG_190; // @[Hold.scala 89:18]
    REG_192 <= REG_191; // @[Hold.scala 89:18]
    REG_193 <= REG_192; // @[Hold.scala 89:18]
    REG_194 <= REG_193; // @[Hold.scala 89:18]
    REG_195 <= REG_194; // @[Hold.scala 89:18]
    REG_196 <= REG_195; // @[Hold.scala 89:18]
    REG_197 <= REG_196; // @[Hold.scala 89:18]
    REG_198 <= REG_197; // @[Hold.scala 89:18]
    REG_199 <= REG_198; // @[Hold.scala 89:18]
    REG_200 <= REG_199; // @[Hold.scala 89:18]
    REG_201 <= REG_200; // @[Hold.scala 89:18]
    REG_202 <= REG_201; // @[Hold.scala 89:18]
    REG_203 <= REG_202; // @[Hold.scala 89:18]
    REG_204 <= REG_203; // @[Hold.scala 89:18]
    REG_205 <= REG_204; // @[Hold.scala 89:18]
    REG_206 <= REG_205; // @[Hold.scala 89:18]
    REG_207 <= REG_206; // @[Hold.scala 89:18]
    REG_208 <= REG_207; // @[Hold.scala 89:18]
    REG_209 <= REG_208; // @[Hold.scala 89:18]
    REG_210 <= REG_209; // @[Hold.scala 89:18]
    REG_211 <= REG_210; // @[Hold.scala 89:18]
    REG_212 <= REG_211; // @[Hold.scala 89:18]
    REG_213 <= REG_212; // @[Hold.scala 89:18]
    REG_214 <= REG_213; // @[Hold.scala 89:18]
    REG_215 <= REG_214; // @[Hold.scala 89:18]
    REG_216 <= REG_215; // @[Hold.scala 89:18]
    REG_217 <= REG_216; // @[Hold.scala 89:18]
    REG_218 <= REG_217; // @[Hold.scala 89:18]
    REG_219 <= REG_218; // @[Hold.scala 89:18]
    REG_220 <= REG_219; // @[Hold.scala 89:18]
    REG_221 <= REG_220; // @[Hold.scala 89:18]
    REG_222 <= REG_221; // @[Hold.scala 89:18]
    REG_223 <= REG_222; // @[Hold.scala 89:18]
    REG_224 <= REG_223; // @[Hold.scala 89:18]
    REG_225 <= REG_224; // @[Hold.scala 89:18]
    REG_226 <= REG_225; // @[Hold.scala 89:18]
    REG_227 <= REG_226; // @[Hold.scala 89:18]
    REG_228 <= REG_227; // @[Hold.scala 89:18]
    REG_229 <= REG_228; // @[Hold.scala 89:18]
    REG_230 <= REG_229; // @[Hold.scala 89:18]
    REG_231 <= REG_230; // @[Hold.scala 89:18]
    REG_232 <= REG_231; // @[Hold.scala 89:18]
    REG_233 <= REG_232; // @[Hold.scala 89:18]
    REG_234 <= REG_233; // @[Hold.scala 89:18]
    REG_235 <= REG_234; // @[Hold.scala 89:18]
    REG_236 <= REG_235; // @[Hold.scala 89:18]
    REG_237 <= REG_236; // @[Hold.scala 89:18]
    REG_238 <= REG_237; // @[Hold.scala 89:18]
    REG_239 <= REG_238; // @[Hold.scala 89:18]
    REG_240 <= REG_239; // @[Hold.scala 89:18]
    REG_241 <= REG_240; // @[Hold.scala 89:18]
    REG_242 <= REG_241; // @[Hold.scala 89:18]
    REG_243 <= REG_242; // @[Hold.scala 89:18]
    REG_244 <= REG_243; // @[Hold.scala 89:18]
    REG_245 <= REG_244; // @[Hold.scala 89:18]
    REG_246 <= REG_245; // @[Hold.scala 89:18]
    REG_247 <= REG_246; // @[Hold.scala 89:18]
    REG_248 <= REG_247; // @[Hold.scala 89:18]
    REG_249 <= REG_248; // @[Hold.scala 89:18]
    REG_250 <= REG_249; // @[Hold.scala 89:18]
    REG_251 <= REG_250; // @[Hold.scala 89:18]
    REG_252 <= REG_251; // @[Hold.scala 89:18]
    REG_253 <= REG_252; // @[Hold.scala 89:18]
    REG_254 <= REG_253; // @[Hold.scala 89:18]
    REG_255 <= REG_254; // @[Hold.scala 89:18]
    REG_256 <= REG_255; // @[Hold.scala 89:18]
    REG_257 <= REG_256; // @[Hold.scala 89:18]
    REG_258 <= REG_257; // @[Hold.scala 89:18]
    REG_259 <= REG_258; // @[Hold.scala 89:18]
    REG_260 <= REG_259; // @[Hold.scala 89:18]
    REG_261 <= REG_260; // @[Hold.scala 89:18]
    REG_262 <= REG_261; // @[Hold.scala 89:18]
    REG_263 <= REG_262; // @[Hold.scala 89:18]
    REG_264 <= REG_263; // @[Hold.scala 89:18]
    REG_265 <= REG_264; // @[Hold.scala 89:18]
    REG_266 <= REG_265; // @[Hold.scala 89:18]
    REG_267 <= REG_266; // @[Hold.scala 89:18]
    REG_268 <= REG_267; // @[Hold.scala 89:18]
    REG_269 <= REG_268; // @[Hold.scala 89:18]
    REG_270 <= REG_269; // @[Hold.scala 89:18]
    REG_271 <= REG_270; // @[Hold.scala 89:18]
    REG_272 <= REG_271; // @[Hold.scala 89:18]
    REG_273 <= REG_272; // @[Hold.scala 89:18]
    REG_274 <= REG_273; // @[Hold.scala 89:18]
    REG_275 <= REG_274; // @[Hold.scala 89:18]
    REG_276 <= REG_275; // @[Hold.scala 89:18]
    REG_277 <= REG_276; // @[Hold.scala 89:18]
    REG_278 <= REG_277; // @[Hold.scala 89:18]
    REG_279 <= REG_278; // @[Hold.scala 89:18]
    REG_280 <= REG_279; // @[Hold.scala 89:18]
    REG_281 <= REG_280; // @[Hold.scala 89:18]
    REG_282 <= REG_281; // @[Hold.scala 89:18]
    REG_283 <= REG_282; // @[Hold.scala 89:18]
    REG_284 <= REG_283; // @[Hold.scala 89:18]
    REG_285 <= REG_284; // @[Hold.scala 89:18]
    REG_286 <= REG_285; // @[Hold.scala 89:18]
    REG_287 <= REG_286; // @[Hold.scala 89:18]
    REG_288 <= REG_287; // @[Hold.scala 89:18]
    REG_289 <= REG_288; // @[Hold.scala 89:18]
    REG_290 <= REG_289; // @[Hold.scala 89:18]
    REG_291 <= REG_290; // @[Hold.scala 89:18]
    REG_292 <= REG_291; // @[Hold.scala 89:18]
    REG_293 <= REG_292; // @[Hold.scala 89:18]
    REG_294 <= REG_293; // @[Hold.scala 89:18]
    REG_295 <= REG_294; // @[Hold.scala 89:18]
    REG_296 <= REG_295; // @[Hold.scala 89:18]
    REG_297 <= REG_296; // @[Hold.scala 89:18]
    REG_298 <= REG_297; // @[Hold.scala 89:18]
    REG_299 <= REG_298; // @[Hold.scala 89:18]
    REG_300 <= REG_299; // @[Hold.scala 89:18]
    REG_301 <= REG_300; // @[Hold.scala 89:18]
    REG_302 <= REG_301; // @[Hold.scala 89:18]
    REG_303 <= REG_302; // @[Hold.scala 89:18]
    REG_304 <= REG_303; // @[Hold.scala 89:18]
    REG_305 <= REG_304; // @[Hold.scala 89:18]
    REG_306 <= REG_305; // @[Hold.scala 89:18]
    REG_307 <= REG_306; // @[Hold.scala 89:18]
    REG_308 <= REG_307; // @[Hold.scala 89:18]
    REG_309 <= REG_308; // @[Hold.scala 89:18]
    REG_310 <= REG_309; // @[Hold.scala 89:18]
    REG_311 <= REG_310; // @[Hold.scala 89:18]
    REG_312 <= REG_311; // @[Hold.scala 89:18]
    REG_313 <= REG_312; // @[Hold.scala 89:18]
    REG_314 <= REG_313; // @[Hold.scala 89:18]
    REG_315 <= REG_314; // @[Hold.scala 89:18]
    REG_316 <= REG_315; // @[Hold.scala 89:18]
    REG_317 <= REG_316; // @[Hold.scala 89:18]
    REG_318 <= REG_317; // @[Hold.scala 89:18]
    REG_319 <= REG_318; // @[Hold.scala 89:18]
    REG_320 <= REG_319; // @[Hold.scala 89:18]
    REG_321 <= REG_320; // @[Hold.scala 89:18]
    REG_322 <= REG_321; // @[Hold.scala 89:18]
    REG_323 <= REG_322; // @[Hold.scala 89:18]
    REG_324 <= REG_323; // @[Hold.scala 89:18]
    REG_325 <= REG_324; // @[Hold.scala 89:18]
    REG_326 <= REG_325; // @[Hold.scala 89:18]
    REG_327 <= REG_326; // @[Hold.scala 89:18]
    REG_328 <= REG_327; // @[Hold.scala 89:18]
    REG_329 <= REG_328; // @[Hold.scala 89:18]
    REG_330 <= REG_329; // @[Hold.scala 89:18]
    REG_331 <= REG_330; // @[Hold.scala 89:18]
    REG_332 <= REG_331; // @[Hold.scala 89:18]
    REG_333 <= REG_332; // @[Hold.scala 89:18]
    REG_334 <= REG_333; // @[Hold.scala 89:18]
    REG_335 <= REG_334; // @[Hold.scala 89:18]
    REG_336 <= REG_335; // @[Hold.scala 89:18]
    REG_337 <= REG_336; // @[Hold.scala 89:18]
    REG_338 <= REG_337; // @[Hold.scala 89:18]
    REG_339 <= REG_338; // @[Hold.scala 89:18]
    REG_340 <= REG_339; // @[Hold.scala 89:18]
    REG_341 <= REG_340; // @[Hold.scala 89:18]
    REG_342 <= REG_341; // @[Hold.scala 89:18]
    REG_343 <= REG_342; // @[Hold.scala 89:18]
    REG_344 <= REG_343; // @[Hold.scala 89:18]
    REG_345 <= REG_344; // @[Hold.scala 89:18]
    REG_346 <= REG_345; // @[Hold.scala 89:18]
    REG_347 <= REG_346; // @[Hold.scala 89:18]
    REG_348 <= REG_347; // @[Hold.scala 89:18]
    REG_349 <= REG_348; // @[Hold.scala 89:18]
    REG_350 <= REG_349; // @[Hold.scala 89:18]
    REG_351 <= REG_350; // @[Hold.scala 89:18]
    REG_352 <= REG_351; // @[Hold.scala 89:18]
    REG_353 <= REG_352; // @[Hold.scala 89:18]
    REG_354 <= REG_353; // @[Hold.scala 89:18]
    REG_355 <= REG_354; // @[Hold.scala 89:18]
    REG_356 <= REG_355; // @[Hold.scala 89:18]
    REG_357 <= REG_356; // @[Hold.scala 89:18]
    REG_358 <= REG_357; // @[Hold.scala 89:18]
    REG_359 <= REG_358; // @[Hold.scala 89:18]
    REG_360 <= REG_359; // @[Hold.scala 89:18]
    REG_361 <= REG_360; // @[Hold.scala 89:18]
    REG_362 <= REG_361; // @[Hold.scala 89:18]
    REG_363 <= REG_362; // @[Hold.scala 89:18]
    REG_364 <= REG_363; // @[Hold.scala 89:18]
    REG_365 <= REG_364; // @[Hold.scala 89:18]
    REG_366 <= REG_365; // @[Hold.scala 89:18]
    REG_367 <= REG_366; // @[Hold.scala 89:18]
    REG_368 <= REG_367; // @[Hold.scala 89:18]
    REG_369 <= REG_368; // @[Hold.scala 89:18]
    REG_370 <= REG_369; // @[Hold.scala 89:18]
    REG_371 <= REG_370; // @[Hold.scala 89:18]
    REG_372 <= REG_371; // @[Hold.scala 89:18]
    REG_373 <= REG_372; // @[Hold.scala 89:18]
    REG_374 <= REG_373; // @[Hold.scala 89:18]
    REG_375 <= REG_374; // @[Hold.scala 89:18]
    REG_376 <= REG_375; // @[Hold.scala 89:18]
    REG_377 <= REG_376; // @[Hold.scala 89:18]
    REG_378 <= REG_377; // @[Hold.scala 89:18]
    REG_379 <= REG_378; // @[Hold.scala 89:18]
    REG_380 <= REG_379; // @[Hold.scala 89:18]
    REG_381 <= REG_380; // @[Hold.scala 89:18]
    REG_382 <= REG_381; // @[Hold.scala 89:18]
    REG_383 <= REG_382; // @[Hold.scala 89:18]
    REG_384 <= REG_383; // @[Hold.scala 89:18]
    REG_385 <= REG_384; // @[Hold.scala 89:18]
    REG_386 <= REG_385; // @[Hold.scala 89:18]
    REG_387 <= REG_386; // @[Hold.scala 89:18]
    REG_388 <= REG_387; // @[Hold.scala 89:18]
    REG_389 <= REG_388; // @[Hold.scala 89:18]
    REG_390 <= REG_389; // @[Hold.scala 89:18]
    REG_391 <= REG_390; // @[Hold.scala 89:18]
    REG_392 <= REG_391; // @[Hold.scala 89:18]
    REG_393 <= REG_392; // @[Hold.scala 89:18]
    REG_394 <= REG_393; // @[Hold.scala 89:18]
    REG_395 <= REG_394; // @[Hold.scala 89:18]
    REG_396 <= REG_395; // @[Hold.scala 89:18]
    REG_397 <= REG_396; // @[Hold.scala 89:18]
    REG_398 <= REG_397; // @[Hold.scala 89:18]
    REG_399 <= REG_398; // @[Hold.scala 89:18]
    REG_400 <= REG_399; // @[Hold.scala 89:18]
    REG_401 <= REG_400; // @[Hold.scala 89:18]
    REG_402 <= REG_401; // @[Hold.scala 89:18]
    REG_403 <= REG_402; // @[Hold.scala 89:18]
    REG_404 <= REG_403; // @[Hold.scala 89:18]
    REG_405 <= REG_404; // @[Hold.scala 89:18]
    REG_406 <= REG_405; // @[Hold.scala 89:18]
    REG_407 <= REG_406; // @[Hold.scala 89:18]
    REG_408 <= REG_407; // @[Hold.scala 89:18]
    REG_409 <= REG_408; // @[Hold.scala 89:18]
    REG_410 <= REG_409; // @[Hold.scala 89:18]
    REG_411 <= REG_410; // @[Hold.scala 89:18]
    REG_412 <= REG_411; // @[Hold.scala 89:18]
    REG_413 <= REG_412; // @[Hold.scala 89:18]
    REG_414 <= REG_413; // @[Hold.scala 89:18]
    REG_415 <= REG_414; // @[Hold.scala 89:18]
    REG_416 <= REG_415; // @[Hold.scala 89:18]
    REG_417 <= REG_416; // @[Hold.scala 89:18]
    REG_418 <= REG_417; // @[Hold.scala 89:18]
    REG_419 <= REG_418; // @[Hold.scala 89:18]
    REG_420 <= REG_419; // @[Hold.scala 89:18]
    REG_421 <= REG_420; // @[Hold.scala 89:18]
    REG_422 <= REG_421; // @[Hold.scala 89:18]
    REG_423 <= REG_422; // @[Hold.scala 89:18]
    REG_424 <= REG_423; // @[Hold.scala 89:18]
    REG_425 <= REG_424; // @[Hold.scala 89:18]
    REG_426 <= REG_425; // @[Hold.scala 89:18]
    REG_427 <= REG_426; // @[Hold.scala 89:18]
    REG_428 <= REG_427; // @[Hold.scala 89:18]
    REG_429 <= REG_428; // @[Hold.scala 89:18]
    REG_430 <= REG_429; // @[Hold.scala 89:18]
    REG_431 <= REG_430; // @[Hold.scala 89:18]
    REG_432 <= REG_431; // @[Hold.scala 89:18]
    REG_433 <= REG_432; // @[Hold.scala 89:18]
    REG_434 <= REG_433; // @[Hold.scala 89:18]
    REG_435 <= REG_434; // @[Hold.scala 89:18]
    REG_436 <= REG_435; // @[Hold.scala 89:18]
    REG_437 <= REG_436; // @[Hold.scala 89:18]
    REG_438 <= REG_437; // @[Hold.scala 89:18]
    REG_439 <= REG_438; // @[Hold.scala 89:18]
    REG_440 <= REG_439; // @[Hold.scala 89:18]
    REG_441 <= REG_440; // @[Hold.scala 89:18]
    REG_442 <= REG_441; // @[Hold.scala 89:18]
    REG_443 <= REG_442; // @[Hold.scala 89:18]
    REG_444 <= REG_443; // @[Hold.scala 89:18]
    REG_445 <= REG_444; // @[Hold.scala 89:18]
    REG_446 <= REG_445; // @[Hold.scala 89:18]
    REG_447 <= REG_446; // @[Hold.scala 89:18]
    REG_448 <= REG_447; // @[Hold.scala 89:18]
    REG_449 <= REG_448; // @[Hold.scala 89:18]
    REG_450 <= REG_449; // @[Hold.scala 89:18]
    REG_451 <= REG_450; // @[Hold.scala 89:18]
    REG_452 <= REG_451; // @[Hold.scala 89:18]
    REG_453 <= REG_452; // @[Hold.scala 89:18]
    REG_454 <= REG_453; // @[Hold.scala 89:18]
    REG_455 <= REG_454; // @[Hold.scala 89:18]
    REG_456 <= REG_455; // @[Hold.scala 89:18]
    REG_457 <= REG_456; // @[Hold.scala 89:18]
    REG_458 <= REG_457; // @[Hold.scala 89:18]
    REG_459 <= REG_458; // @[Hold.scala 89:18]
    REG_460 <= REG_459; // @[Hold.scala 89:18]
    REG_461 <= REG_460; // @[Hold.scala 89:18]
    REG_462 <= REG_461; // @[Hold.scala 89:18]
    REG_463 <= REG_462; // @[Hold.scala 89:18]
    REG_464 <= REG_463; // @[Hold.scala 89:18]
    REG_465 <= REG_464; // @[Hold.scala 89:18]
    REG_466 <= REG_465; // @[Hold.scala 89:18]
    REG_467 <= REG_466; // @[Hold.scala 89:18]
    REG_468 <= REG_467; // @[Hold.scala 89:18]
    REG_469 <= REG_468; // @[Hold.scala 89:18]
    REG_470 <= REG_469; // @[Hold.scala 89:18]
    REG_471 <= REG_470; // @[Hold.scala 89:18]
    REG_472 <= REG_471; // @[Hold.scala 89:18]
    REG_473 <= REG_472; // @[Hold.scala 89:18]
    REG_474 <= REG_473; // @[Hold.scala 89:18]
    REG_475 <= REG_474; // @[Hold.scala 89:18]
    REG_476 <= REG_475; // @[Hold.scala 89:18]
    REG_477 <= REG_476; // @[Hold.scala 89:18]
    REG_478 <= REG_477; // @[Hold.scala 89:18]
    REG_479 <= REG_478; // @[Hold.scala 89:18]
    REG_480 <= REG_479; // @[Hold.scala 89:18]
    REG_481 <= REG_480; // @[Hold.scala 89:18]
    REG_482 <= REG_481; // @[Hold.scala 89:18]
    REG_483 <= REG_482; // @[Hold.scala 89:18]
    REG_484 <= REG_483; // @[Hold.scala 89:18]
    REG_485 <= REG_484; // @[Hold.scala 89:18]
    REG_486 <= REG_485; // @[Hold.scala 89:18]
    REG_487 <= REG_486; // @[Hold.scala 89:18]
    REG_488 <= REG_487; // @[Hold.scala 89:18]
    REG_489 <= REG_488; // @[Hold.scala 89:18]
    REG_490 <= REG_489; // @[Hold.scala 89:18]
    REG_491 <= REG_490; // @[Hold.scala 89:18]
    REG_492 <= REG_491; // @[Hold.scala 89:18]
    REG_493 <= REG_492; // @[Hold.scala 89:18]
    REG_494 <= REG_493; // @[Hold.scala 89:18]
    REG_495 <= REG_494; // @[Hold.scala 89:18]
    REG_496 <= REG_495; // @[Hold.scala 89:18]
    REG_497 <= REG_496; // @[Hold.scala 89:18]
    REG_498 <= REG_497; // @[Hold.scala 89:18]
    REG_499 <= REG_498; // @[Hold.scala 89:18]
    REG_500 <= REG_499; // @[Hold.scala 89:18]
    REG_501 <= REG_500; // @[Hold.scala 89:18]
    REG_502 <= REG_501; // @[Hold.scala 89:18]
    REG_503 <= REG_502; // @[Hold.scala 89:18]
    REG_504 <= REG_503; // @[Hold.scala 89:18]
    REG_505 <= REG_504; // @[Hold.scala 89:18]
    REG_506 <= REG_505; // @[Hold.scala 89:18]
    REG_507 <= REG_506; // @[Hold.scala 89:18]
    REG_508 <= REG_507; // @[Hold.scala 89:18]
    REG_509 <= REG_508; // @[Hold.scala 89:18]
    REG_510 <= REG_509; // @[Hold.scala 89:18]
    REG_511 <= REG_510; // @[Hold.scala 89:18]
    REG_512 <= REG_511; // @[Hold.scala 89:18]
    REG_513 <= REG_512; // @[Hold.scala 89:18]
    REG_514 <= REG_513; // @[Hold.scala 89:18]
    REG_515 <= REG_514; // @[Hold.scala 89:18]
    REG_516 <= REG_515; // @[Hold.scala 89:18]
    REG_517 <= REG_516; // @[Hold.scala 89:18]
    REG_518 <= REG_517; // @[Hold.scala 89:18]
    REG_519 <= REG_518; // @[Hold.scala 89:18]
    REG_520 <= REG_519; // @[Hold.scala 89:18]
    REG_521 <= REG_520; // @[Hold.scala 89:18]
    REG_522 <= REG_521; // @[Hold.scala 89:18]
    REG_523 <= REG_522; // @[Hold.scala 89:18]
    REG_524 <= REG_523; // @[Hold.scala 89:18]
    REG_525 <= REG_524; // @[Hold.scala 89:18]
    REG_526 <= REG_525; // @[Hold.scala 89:18]
    REG_527 <= REG_526; // @[Hold.scala 89:18]
    REG_528 <= REG_527; // @[Hold.scala 89:18]
    REG_529 <= REG_528; // @[Hold.scala 89:18]
    REG_530 <= REG_529; // @[Hold.scala 89:18]
    REG_531 <= REG_530; // @[Hold.scala 89:18]
    REG_532 <= REG_531; // @[Hold.scala 89:18]
    REG_533 <= REG_532; // @[Hold.scala 89:18]
    REG_534 <= REG_533; // @[Hold.scala 89:18]
    REG_535 <= REG_534; // @[Hold.scala 89:18]
    REG_536 <= REG_535; // @[Hold.scala 89:18]
    REG_537 <= REG_536; // @[Hold.scala 89:18]
    REG_538 <= REG_537; // @[Hold.scala 89:18]
    REG_539 <= REG_538; // @[Hold.scala 89:18]
    REG_540 <= REG_539; // @[Hold.scala 89:18]
    REG_541 <= REG_540; // @[Hold.scala 89:18]
    REG_542 <= REG_541; // @[Hold.scala 89:18]
    REG_543 <= REG_542; // @[Hold.scala 89:18]
    REG_544 <= REG_543; // @[Hold.scala 89:18]
    REG_545 <= REG_544; // @[Hold.scala 89:18]
    REG_546 <= REG_545; // @[Hold.scala 89:18]
    REG_547 <= REG_546; // @[Hold.scala 89:18]
    REG_548 <= REG_547; // @[Hold.scala 89:18]
    REG_549 <= REG_548; // @[Hold.scala 89:18]
    REG_550 <= REG_549; // @[Hold.scala 89:18]
    REG_551 <= REG_550; // @[Hold.scala 89:18]
    REG_552 <= REG_551; // @[Hold.scala 89:18]
    REG_553 <= REG_552; // @[Hold.scala 89:18]
    REG_554 <= REG_553; // @[Hold.scala 89:18]
    REG_555 <= REG_554; // @[Hold.scala 89:18]
    REG_556 <= REG_555; // @[Hold.scala 89:18]
    REG_557 <= REG_556; // @[Hold.scala 89:18]
    REG_558 <= REG_557; // @[Hold.scala 89:18]
    REG_559 <= REG_558; // @[Hold.scala 89:18]
    REG_560 <= REG_559; // @[Hold.scala 89:18]
    REG_561 <= REG_560; // @[Hold.scala 89:18]
    REG_562 <= REG_561; // @[Hold.scala 89:18]
    REG_563 <= REG_562; // @[Hold.scala 89:18]
    REG_564 <= REG_563; // @[Hold.scala 89:18]
    REG_565 <= REG_564; // @[Hold.scala 89:18]
    REG_566 <= REG_565; // @[Hold.scala 89:18]
    REG_567 <= REG_566; // @[Hold.scala 89:18]
    REG_568 <= REG_567; // @[Hold.scala 89:18]
    REG_569 <= REG_568; // @[Hold.scala 89:18]
    REG_570 <= REG_569; // @[Hold.scala 89:18]
    REG_571 <= REG_570; // @[Hold.scala 89:18]
    REG_572 <= REG_571; // @[Hold.scala 89:18]
    REG_573 <= REG_572; // @[Hold.scala 89:18]
    REG_574 <= REG_573; // @[Hold.scala 89:18]
    REG_575 <= REG_574; // @[Hold.scala 89:18]
    REG_576 <= REG_575; // @[Hold.scala 89:18]
    REG_577 <= REG_576; // @[Hold.scala 89:18]
    REG_578 <= REG_577; // @[Hold.scala 89:18]
    REG_579 <= REG_578; // @[Hold.scala 89:18]
    REG_580 <= REG_579; // @[Hold.scala 89:18]
    REG_581 <= REG_580; // @[Hold.scala 89:18]
    REG_582 <= REG_581; // @[Hold.scala 89:18]
    REG_583 <= REG_582; // @[Hold.scala 89:18]
    REG_584 <= REG_583; // @[Hold.scala 89:18]
    REG_585 <= REG_584; // @[Hold.scala 89:18]
    REG_586 <= REG_585; // @[Hold.scala 89:18]
    REG_587 <= REG_586; // @[Hold.scala 89:18]
    REG_588 <= REG_587; // @[Hold.scala 89:18]
    REG_589 <= REG_588; // @[Hold.scala 89:18]
    REG_590 <= REG_589; // @[Hold.scala 89:18]
    REG_591 <= REG_590; // @[Hold.scala 89:18]
    REG_592 <= REG_591; // @[Hold.scala 89:18]
    REG_593 <= REG_592; // @[Hold.scala 89:18]
    REG_594 <= REG_593; // @[Hold.scala 89:18]
    REG_595 <= REG_594; // @[Hold.scala 89:18]
    REG_596 <= REG_595; // @[Hold.scala 89:18]
    REG_597 <= REG_596; // @[Hold.scala 89:18]
    REG_598 <= REG_597; // @[Hold.scala 89:18]
    REG_599 <= REG_598; // @[Hold.scala 89:18]
    REG_600 <= REG_599; // @[Hold.scala 89:18]
    REG_601 <= REG_600; // @[Hold.scala 89:18]
    REG_602 <= REG_601; // @[Hold.scala 89:18]
    REG_603 <= REG_602; // @[Hold.scala 89:18]
    REG_604 <= REG_603; // @[Hold.scala 89:18]
    REG_605 <= REG_604; // @[Hold.scala 89:18]
    REG_606 <= REG_605; // @[Hold.scala 89:18]
    REG_607 <= REG_606; // @[Hold.scala 89:18]
    REG_608 <= REG_607; // @[Hold.scala 89:18]
    REG_609 <= REG_608; // @[Hold.scala 89:18]
    REG_610 <= REG_609; // @[Hold.scala 89:18]
    REG_611 <= REG_610; // @[Hold.scala 89:18]
    REG_612 <= REG_611; // @[Hold.scala 89:18]
    REG_613 <= REG_612; // @[Hold.scala 89:18]
    REG_614 <= REG_613; // @[Hold.scala 89:18]
    REG_615 <= REG_614; // @[Hold.scala 89:18]
    REG_616 <= REG_615; // @[Hold.scala 89:18]
    REG_617 <= REG_616; // @[Hold.scala 89:18]
    REG_618 <= REG_617; // @[Hold.scala 89:18]
    REG_619 <= REG_618; // @[Hold.scala 89:18]
    REG_620 <= REG_619; // @[Hold.scala 89:18]
    REG_621 <= REG_620; // @[Hold.scala 89:18]
    REG_622 <= REG_621; // @[Hold.scala 89:18]
    REG_623 <= REG_622; // @[Hold.scala 89:18]
    REG_624 <= REG_623; // @[Hold.scala 89:18]
    REG_625 <= REG_624; // @[Hold.scala 89:18]
    REG_626 <= REG_625; // @[Hold.scala 89:18]
    REG_627 <= REG_626; // @[Hold.scala 89:18]
    REG_628 <= REG_627; // @[Hold.scala 89:18]
    REG_629 <= REG_628; // @[Hold.scala 89:18]
    REG_630 <= REG_629; // @[Hold.scala 89:18]
    REG_631 <= REG_630; // @[Hold.scala 89:18]
    REG_632 <= REG_631; // @[Hold.scala 89:18]
    REG_633 <= REG_632; // @[Hold.scala 89:18]
    REG_634 <= REG_633; // @[Hold.scala 89:18]
    REG_635 <= REG_634; // @[Hold.scala 89:18]
    REG_636 <= REG_635; // @[Hold.scala 89:18]
    REG_637 <= REG_636; // @[Hold.scala 89:18]
    REG_638 <= REG_637; // @[Hold.scala 89:18]
    REG_639 <= REG_638; // @[Hold.scala 89:18]
    REG_640 <= REG_639; // @[Hold.scala 89:18]
    REG_641 <= REG_640; // @[Hold.scala 89:18]
    REG_642 <= REG_641; // @[Hold.scala 89:18]
    REG_643 <= REG_642; // @[Hold.scala 89:18]
    REG_644 <= REG_643; // @[Hold.scala 89:18]
    REG_645 <= REG_644; // @[Hold.scala 89:18]
    REG_646 <= REG_645; // @[Hold.scala 89:18]
    REG_647 <= REG_646; // @[Hold.scala 89:18]
    REG_648 <= REG_647; // @[Hold.scala 89:18]
    REG_649 <= REG_648; // @[Hold.scala 89:18]
    REG_650 <= REG_649; // @[Hold.scala 89:18]
    REG_651 <= REG_650; // @[Hold.scala 89:18]
    REG_652 <= REG_651; // @[Hold.scala 89:18]
    REG_653 <= REG_652; // @[Hold.scala 89:18]
    REG_654 <= REG_653; // @[Hold.scala 89:18]
    REG_655 <= REG_654; // @[Hold.scala 89:18]
    REG_656 <= REG_655; // @[Hold.scala 89:18]
    REG_657 <= REG_656; // @[Hold.scala 89:18]
    REG_658 <= REG_657; // @[Hold.scala 89:18]
    REG_659 <= REG_658; // @[Hold.scala 89:18]
    REG_660 <= REG_659; // @[Hold.scala 89:18]
    REG_661 <= REG_660; // @[Hold.scala 89:18]
    REG_662 <= REG_661; // @[Hold.scala 89:18]
    REG_663 <= REG_662; // @[Hold.scala 89:18]
    REG_664 <= REG_663; // @[Hold.scala 89:18]
    REG_665 <= REG_664; // @[Hold.scala 89:18]
    REG_666 <= REG_665; // @[Hold.scala 89:18]
    REG_667 <= REG_666; // @[Hold.scala 89:18]
    REG_668 <= REG_667; // @[Hold.scala 89:18]
    REG_669 <= REG_668; // @[Hold.scala 89:18]
    REG_670 <= REG_669; // @[Hold.scala 89:18]
    REG_671 <= REG_670; // @[Hold.scala 89:18]
    REG_672 <= REG_671; // @[Hold.scala 89:18]
    REG_673 <= REG_672; // @[Hold.scala 89:18]
    REG_674 <= REG_673; // @[Hold.scala 89:18]
    REG_675 <= REG_674; // @[Hold.scala 89:18]
    REG_676 <= REG_675; // @[Hold.scala 89:18]
    REG_677 <= REG_676; // @[Hold.scala 89:18]
    REG_678 <= REG_677; // @[Hold.scala 89:18]
    REG_679 <= REG_678; // @[Hold.scala 89:18]
    REG_680 <= REG_679; // @[Hold.scala 89:18]
    REG_681 <= REG_680; // @[Hold.scala 89:18]
    REG_682 <= REG_681; // @[Hold.scala 89:18]
    REG_683 <= REG_682; // @[Hold.scala 89:18]
    REG_684 <= REG_683; // @[Hold.scala 89:18]
    REG_685 <= REG_684; // @[Hold.scala 89:18]
    REG_686 <= REG_685; // @[Hold.scala 89:18]
    REG_687 <= REG_686; // @[Hold.scala 89:18]
    REG_688 <= REG_687; // @[Hold.scala 89:18]
    REG_689 <= REG_688; // @[Hold.scala 89:18]
    REG_690 <= REG_689; // @[Hold.scala 89:18]
    REG_691 <= REG_690; // @[Hold.scala 89:18]
    REG_692 <= REG_691; // @[Hold.scala 89:18]
    REG_693 <= REG_692; // @[Hold.scala 89:18]
    REG_694 <= REG_693; // @[Hold.scala 89:18]
    REG_695 <= REG_694; // @[Hold.scala 89:18]
    REG_696 <= REG_695; // @[Hold.scala 89:18]
    REG_697 <= REG_696; // @[Hold.scala 89:18]
    REG_698 <= REG_697; // @[Hold.scala 89:18]
    REG_699 <= REG_698; // @[Hold.scala 89:18]
    REG_700 <= REG_699; // @[Hold.scala 89:18]
    REG_701 <= REG_700; // @[Hold.scala 89:18]
    REG_702 <= REG_701; // @[Hold.scala 89:18]
    REG_703 <= REG_702; // @[Hold.scala 89:18]
    REG_704 <= REG_703; // @[Hold.scala 89:18]
    REG_705 <= REG_704; // @[Hold.scala 89:18]
    REG_706 <= REG_705; // @[Hold.scala 89:18]
    REG_707 <= REG_706; // @[Hold.scala 89:18]
    REG_708 <= REG_707; // @[Hold.scala 89:18]
    REG_709 <= REG_708; // @[Hold.scala 89:18]
    REG_710 <= REG_709; // @[Hold.scala 89:18]
    REG_711 <= REG_710; // @[Hold.scala 89:18]
    REG_712 <= REG_711; // @[Hold.scala 89:18]
    REG_713 <= REG_712; // @[Hold.scala 89:18]
    REG_714 <= REG_713; // @[Hold.scala 89:18]
    REG_715 <= REG_714; // @[Hold.scala 89:18]
    REG_716 <= REG_715; // @[Hold.scala 89:18]
    REG_717 <= REG_716; // @[Hold.scala 89:18]
    REG_718 <= REG_717; // @[Hold.scala 89:18]
    REG_719 <= REG_718; // @[Hold.scala 89:18]
    REG_720 <= REG_719; // @[Hold.scala 89:18]
    REG_721 <= REG_720; // @[Hold.scala 89:18]
    REG_722 <= REG_721; // @[Hold.scala 89:18]
    REG_723 <= REG_722; // @[Hold.scala 89:18]
    REG_724 <= REG_723; // @[Hold.scala 89:18]
    REG_725 <= REG_724; // @[Hold.scala 89:18]
    REG_726 <= REG_725; // @[Hold.scala 89:18]
    REG_727 <= REG_726; // @[Hold.scala 89:18]
    REG_728 <= REG_727; // @[Hold.scala 89:18]
    REG_729 <= REG_728; // @[Hold.scala 89:18]
    REG_730 <= REG_729; // @[Hold.scala 89:18]
    REG_731 <= REG_730; // @[Hold.scala 89:18]
    REG_732 <= REG_731; // @[Hold.scala 89:18]
    REG_733 <= REG_732; // @[Hold.scala 89:18]
    REG_734 <= REG_733; // @[Hold.scala 89:18]
    REG_735 <= REG_734; // @[Hold.scala 89:18]
    REG_736 <= REG_735; // @[Hold.scala 89:18]
    REG_737 <= REG_736; // @[Hold.scala 89:18]
    REG_738 <= REG_737; // @[Hold.scala 89:18]
    REG_739 <= REG_738; // @[Hold.scala 89:18]
    REG_740 <= REG_739; // @[Hold.scala 89:18]
    REG_741 <= REG_740; // @[Hold.scala 89:18]
    REG_742 <= REG_741; // @[Hold.scala 89:18]
    REG_743 <= REG_742; // @[Hold.scala 89:18]
    REG_744 <= REG_743; // @[Hold.scala 89:18]
    REG_745 <= REG_744; // @[Hold.scala 89:18]
    REG_746 <= REG_745; // @[Hold.scala 89:18]
    REG_747 <= REG_746; // @[Hold.scala 89:18]
    REG_748 <= REG_747; // @[Hold.scala 89:18]
    REG_749 <= REG_748; // @[Hold.scala 89:18]
    REG_750 <= REG_749; // @[Hold.scala 89:18]
    REG_751 <= REG_750; // @[Hold.scala 89:18]
    REG_752 <= REG_751; // @[Hold.scala 89:18]
    REG_753 <= REG_752; // @[Hold.scala 89:18]
    REG_754 <= REG_753; // @[Hold.scala 89:18]
    REG_755 <= REG_754; // @[Hold.scala 89:18]
    REG_756 <= REG_755; // @[Hold.scala 89:18]
    REG_757 <= REG_756; // @[Hold.scala 89:18]
    REG_758 <= REG_757; // @[Hold.scala 89:18]
    REG_759 <= REG_758; // @[Hold.scala 89:18]
    REG_760 <= REG_759; // @[Hold.scala 89:18]
    REG_761 <= REG_760; // @[Hold.scala 89:18]
    REG_762 <= REG_761; // @[Hold.scala 89:18]
    REG_763 <= REG_762; // @[Hold.scala 89:18]
    REG_764 <= REG_763; // @[Hold.scala 89:18]
    REG_765 <= REG_764; // @[Hold.scala 89:18]
    REG_766 <= REG_765; // @[Hold.scala 89:18]
    REG_767 <= REG_766; // @[Hold.scala 89:18]
    REG_768 <= REG_767; // @[Hold.scala 89:18]
    REG_769 <= REG_768; // @[Hold.scala 89:18]
    REG_770 <= REG_769; // @[Hold.scala 89:18]
    REG_771 <= REG_770; // @[Hold.scala 89:18]
    REG_772 <= REG_771; // @[Hold.scala 89:18]
    REG_773 <= REG_772; // @[Hold.scala 89:18]
    REG_774 <= REG_773; // @[Hold.scala 89:18]
    REG_775 <= REG_774; // @[Hold.scala 89:18]
    REG_776 <= REG_775; // @[Hold.scala 89:18]
    REG_777 <= REG_776; // @[Hold.scala 89:18]
    REG_778 <= REG_777; // @[Hold.scala 89:18]
    REG_779 <= REG_778; // @[Hold.scala 89:18]
    REG_780 <= REG_779; // @[Hold.scala 89:18]
    REG_781 <= REG_780; // @[Hold.scala 89:18]
    REG_782 <= REG_781; // @[Hold.scala 89:18]
    REG_783 <= REG_782; // @[Hold.scala 89:18]
    REG_784 <= REG_783; // @[Hold.scala 89:18]
    REG_785 <= REG_784; // @[Hold.scala 89:18]
    REG_786 <= REG_785; // @[Hold.scala 89:18]
    REG_787 <= REG_786; // @[Hold.scala 89:18]
    REG_788 <= REG_787; // @[Hold.scala 89:18]
    REG_789 <= REG_788; // @[Hold.scala 89:18]
    REG_790 <= REG_789; // @[Hold.scala 89:18]
    REG_791 <= REG_790; // @[Hold.scala 89:18]
    REG_792 <= REG_791; // @[Hold.scala 89:18]
    REG_793 <= REG_792; // @[Hold.scala 89:18]
    REG_794 <= REG_793; // @[Hold.scala 89:18]
    REG_795 <= REG_794; // @[Hold.scala 89:18]
    REG_796 <= REG_795; // @[Hold.scala 89:18]
    REG_797 <= REG_796; // @[Hold.scala 89:18]
    REG_798 <= REG_797; // @[Hold.scala 89:18]
    REG_799 <= REG_798; // @[Hold.scala 89:18]
    REG_800 <= REG_799; // @[Hold.scala 89:18]
    REG_801 <= REG_800; // @[Hold.scala 89:18]
    REG_802 <= REG_801; // @[Hold.scala 89:18]
    REG_803 <= REG_802; // @[Hold.scala 89:18]
    REG_804 <= REG_803; // @[Hold.scala 89:18]
    REG_805 <= REG_804; // @[Hold.scala 89:18]
    REG_806 <= REG_805; // @[Hold.scala 89:18]
    REG_807 <= REG_806; // @[Hold.scala 89:18]
    REG_808 <= REG_807; // @[Hold.scala 89:18]
    REG_809 <= REG_808; // @[Hold.scala 89:18]
    REG_810 <= REG_809; // @[Hold.scala 89:18]
    REG_811 <= REG_810; // @[Hold.scala 89:18]
    REG_812 <= REG_811; // @[Hold.scala 89:18]
    REG_813 <= REG_812; // @[Hold.scala 89:18]
    REG_814 <= REG_813; // @[Hold.scala 89:18]
    REG_815 <= REG_814; // @[Hold.scala 89:18]
    REG_816 <= REG_815; // @[Hold.scala 89:18]
    REG_817 <= REG_816; // @[Hold.scala 89:18]
    REG_818 <= REG_817; // @[Hold.scala 89:18]
    REG_819 <= REG_818; // @[Hold.scala 89:18]
    REG_820 <= REG_819; // @[Hold.scala 89:18]
    REG_821 <= REG_820; // @[Hold.scala 89:18]
    REG_822 <= REG_821; // @[Hold.scala 89:18]
    REG_823 <= REG_822; // @[Hold.scala 89:18]
    REG_824 <= REG_823; // @[Hold.scala 89:18]
    REG_825 <= REG_824; // @[Hold.scala 89:18]
    REG_826 <= REG_825; // @[Hold.scala 89:18]
    REG_827 <= REG_826; // @[Hold.scala 89:18]
    REG_828 <= REG_827; // @[Hold.scala 89:18]
    REG_829 <= REG_828; // @[Hold.scala 89:18]
    REG_830 <= REG_829; // @[Hold.scala 89:18]
    REG_831 <= REG_830; // @[Hold.scala 89:18]
    REG_832 <= REG_831; // @[Hold.scala 89:18]
    REG_833 <= REG_832; // @[Hold.scala 89:18]
    REG_834 <= REG_833; // @[Hold.scala 89:18]
    REG_835 <= REG_834; // @[Hold.scala 89:18]
    REG_836 <= REG_835; // @[Hold.scala 89:18]
    REG_837 <= REG_836; // @[Hold.scala 89:18]
    REG_838 <= REG_837; // @[Hold.scala 89:18]
    REG_839 <= REG_838; // @[Hold.scala 89:18]
    REG_840 <= REG_839; // @[Hold.scala 89:18]
    REG_841 <= REG_840; // @[Hold.scala 89:18]
    REG_842 <= REG_841; // @[Hold.scala 89:18]
    REG_843 <= REG_842; // @[Hold.scala 89:18]
    REG_844 <= REG_843; // @[Hold.scala 89:18]
    REG_845 <= REG_844; // @[Hold.scala 89:18]
    REG_846 <= REG_845; // @[Hold.scala 89:18]
    REG_847 <= REG_846; // @[Hold.scala 89:18]
    REG_848 <= REG_847; // @[Hold.scala 89:18]
    REG_849 <= REG_848; // @[Hold.scala 89:18]
    REG_850 <= REG_849; // @[Hold.scala 89:18]
    REG_851 <= REG_850; // @[Hold.scala 89:18]
    REG_852 <= REG_851; // @[Hold.scala 89:18]
    REG_853 <= REG_852; // @[Hold.scala 89:18]
    REG_854 <= REG_853; // @[Hold.scala 89:18]
    REG_855 <= REG_854; // @[Hold.scala 89:18]
    REG_856 <= REG_855; // @[Hold.scala 89:18]
    REG_857 <= REG_856; // @[Hold.scala 89:18]
    REG_858 <= REG_857; // @[Hold.scala 89:18]
    REG_859 <= REG_858; // @[Hold.scala 89:18]
    REG_860 <= REG_859; // @[Hold.scala 89:18]
    REG_861 <= REG_860; // @[Hold.scala 89:18]
    REG_862 <= REG_861; // @[Hold.scala 89:18]
    REG_863 <= REG_862; // @[Hold.scala 89:18]
    REG_864 <= REG_863; // @[Hold.scala 89:18]
    REG_865 <= REG_864; // @[Hold.scala 89:18]
    REG_866 <= REG_865; // @[Hold.scala 89:18]
    REG_867 <= REG_866; // @[Hold.scala 89:18]
    REG_868 <= REG_867; // @[Hold.scala 89:18]
    REG_869 <= REG_868; // @[Hold.scala 89:18]
    REG_870 <= REG_869; // @[Hold.scala 89:18]
    REG_871 <= REG_870; // @[Hold.scala 89:18]
    REG_872 <= REG_871; // @[Hold.scala 89:18]
    REG_873 <= REG_872; // @[Hold.scala 89:18]
    REG_874 <= REG_873; // @[Hold.scala 89:18]
    REG_875 <= REG_874; // @[Hold.scala 89:18]
    REG_876 <= REG_875; // @[Hold.scala 89:18]
    REG_877 <= REG_876; // @[Hold.scala 89:18]
    REG_878 <= REG_877; // @[Hold.scala 89:18]
    REG_879 <= REG_878; // @[Hold.scala 89:18]
    REG_880 <= REG_879; // @[Hold.scala 89:18]
    REG_881 <= REG_880; // @[Hold.scala 89:18]
    REG_882 <= REG_881; // @[Hold.scala 89:18]
    REG_883 <= REG_882; // @[Hold.scala 89:18]
    REG_884 <= REG_883; // @[Hold.scala 89:18]
    REG_885 <= REG_884; // @[Hold.scala 89:18]
    REG_886 <= REG_885; // @[Hold.scala 89:18]
    REG_887 <= REG_886; // @[Hold.scala 89:18]
    REG_888 <= REG_887; // @[Hold.scala 89:18]
    REG_889 <= REG_888; // @[Hold.scala 89:18]
    REG_890 <= REG_889; // @[Hold.scala 89:18]
    REG_891 <= REG_890; // @[Hold.scala 89:18]
    REG_892 <= REG_891; // @[Hold.scala 89:18]
    REG_893 <= REG_892; // @[Hold.scala 89:18]
    REG_894 <= REG_893; // @[Hold.scala 89:18]
    REG_895 <= REG_894; // @[Hold.scala 89:18]
    REG_896 <= REG_895; // @[Hold.scala 89:18]
    REG_897 <= REG_896; // @[Hold.scala 89:18]
    REG_898 <= REG_897; // @[Hold.scala 89:18]
    REG_899 <= REG_898; // @[Hold.scala 89:18]
    REG_900 <= REG_899; // @[Hold.scala 89:18]
    REG_901 <= REG_900; // @[Hold.scala 89:18]
    REG_902 <= REG_901; // @[Hold.scala 89:18]
    REG_903 <= REG_902; // @[Hold.scala 89:18]
    REG_904 <= REG_903; // @[Hold.scala 89:18]
    REG_905 <= REG_904; // @[Hold.scala 89:18]
    REG_906 <= REG_905; // @[Hold.scala 89:18]
    REG_907 <= REG_906; // @[Hold.scala 89:18]
    REG_908 <= REG_907; // @[Hold.scala 89:18]
    REG_909 <= REG_908; // @[Hold.scala 89:18]
    REG_910 <= REG_909; // @[Hold.scala 89:18]
    REG_911 <= REG_910; // @[Hold.scala 89:18]
    REG_912 <= REG_911; // @[Hold.scala 89:18]
    REG_913 <= REG_912; // @[Hold.scala 89:18]
    REG_914 <= REG_913; // @[Hold.scala 89:18]
    REG_915 <= REG_914; // @[Hold.scala 89:18]
    REG_916 <= REG_915; // @[Hold.scala 89:18]
    REG_917 <= REG_916; // @[Hold.scala 89:18]
    REG_918 <= REG_917; // @[Hold.scala 89:18]
    REG_919 <= REG_918; // @[Hold.scala 89:18]
    REG_920 <= REG_919; // @[Hold.scala 89:18]
    REG_921 <= REG_920; // @[Hold.scala 89:18]
    REG_922 <= REG_921; // @[Hold.scala 89:18]
    REG_923 <= REG_922; // @[Hold.scala 89:18]
    REG_924 <= REG_923; // @[Hold.scala 89:18]
    REG_925 <= REG_924; // @[Hold.scala 89:18]
    REG_926 <= REG_925; // @[Hold.scala 89:18]
    REG_927 <= REG_926; // @[Hold.scala 89:18]
    REG_928 <= REG_927; // @[Hold.scala 89:18]
    REG_929 <= REG_928; // @[Hold.scala 89:18]
    REG_930 <= REG_929; // @[Hold.scala 89:18]
    REG_931 <= REG_930; // @[Hold.scala 89:18]
    REG_932 <= REG_931; // @[Hold.scala 89:18]
    REG_933 <= REG_932; // @[Hold.scala 89:18]
    REG_934 <= REG_933; // @[Hold.scala 89:18]
    REG_935 <= REG_934; // @[Hold.scala 89:18]
    REG_936 <= REG_935; // @[Hold.scala 89:18]
    REG_937 <= REG_936; // @[Hold.scala 89:18]
    REG_938 <= REG_937; // @[Hold.scala 89:18]
    REG_939 <= REG_938; // @[Hold.scala 89:18]
    REG_940 <= REG_939; // @[Hold.scala 89:18]
    REG_941 <= REG_940; // @[Hold.scala 89:18]
    REG_942 <= REG_941; // @[Hold.scala 89:18]
    REG_943 <= REG_942; // @[Hold.scala 89:18]
    REG_944 <= REG_943; // @[Hold.scala 89:18]
    REG_945 <= REG_944; // @[Hold.scala 89:18]
    REG_946 <= REG_945; // @[Hold.scala 89:18]
    REG_947 <= REG_946; // @[Hold.scala 89:18]
    REG_948 <= REG_947; // @[Hold.scala 89:18]
    REG_949 <= REG_948; // @[Hold.scala 89:18]
    REG_950 <= REG_949; // @[Hold.scala 89:18]
    REG_951 <= REG_950; // @[Hold.scala 89:18]
    REG_952 <= REG_951; // @[Hold.scala 89:18]
    REG_953 <= REG_952; // @[Hold.scala 89:18]
    REG_954 <= REG_953; // @[Hold.scala 89:18]
    REG_955 <= REG_954; // @[Hold.scala 89:18]
    REG_956 <= REG_955; // @[Hold.scala 89:18]
    REG_957 <= REG_956; // @[Hold.scala 89:18]
    REG_958 <= REG_957; // @[Hold.scala 89:18]
    REG_959 <= REG_958; // @[Hold.scala 89:18]
    REG_960 <= REG_959; // @[Hold.scala 89:18]
    REG_961 <= REG_960; // @[Hold.scala 89:18]
    REG_962 <= REG_961; // @[Hold.scala 89:18]
    REG_963 <= REG_962; // @[Hold.scala 89:18]
    REG_964 <= REG_963; // @[Hold.scala 89:18]
    REG_965 <= REG_964; // @[Hold.scala 89:18]
    REG_966 <= REG_965; // @[Hold.scala 89:18]
    REG_967 <= REG_966; // @[Hold.scala 89:18]
    REG_968 <= REG_967; // @[Hold.scala 89:18]
    REG_969 <= REG_968; // @[Hold.scala 89:18]
    REG_970 <= REG_969; // @[Hold.scala 89:18]
    REG_971 <= REG_970; // @[Hold.scala 89:18]
    REG_972 <= REG_971; // @[Hold.scala 89:18]
    REG_973 <= REG_972; // @[Hold.scala 89:18]
    REG_974 <= REG_973; // @[Hold.scala 89:18]
    REG_975 <= REG_974; // @[Hold.scala 89:18]
    REG_976 <= REG_975; // @[Hold.scala 89:18]
    REG_977 <= REG_976; // @[Hold.scala 89:18]
    REG_978 <= REG_977; // @[Hold.scala 89:18]
    REG_979 <= REG_978; // @[Hold.scala 89:18]
    REG_980 <= REG_979; // @[Hold.scala 89:18]
    REG_981 <= REG_980; // @[Hold.scala 89:18]
    REG_982 <= REG_981; // @[Hold.scala 89:18]
    REG_983 <= REG_982; // @[Hold.scala 89:18]
    REG_984 <= REG_983; // @[Hold.scala 89:18]
    REG_985 <= REG_984; // @[Hold.scala 89:18]
    REG_986 <= REG_985; // @[Hold.scala 89:18]
    REG_987 <= REG_986; // @[Hold.scala 89:18]
    REG_988 <= REG_987; // @[Hold.scala 89:18]
    REG_989 <= REG_988; // @[Hold.scala 89:18]
    REG_990 <= REG_989; // @[Hold.scala 89:18]
    REG_991 <= REG_990; // @[Hold.scala 89:18]
    REG_992 <= REG_991; // @[Hold.scala 89:18]
    REG_993 <= REG_992; // @[Hold.scala 89:18]
    REG_994 <= REG_993; // @[Hold.scala 89:18]
    REG_995 <= REG_994; // @[Hold.scala 89:18]
    REG_996 <= REG_995; // @[Hold.scala 89:18]
    REG_997 <= REG_996; // @[Hold.scala 89:18]
    REG_998 <= REG_997; // @[Hold.scala 89:18]
    out <= REG_998; // @[Hold.scala 89:18]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  REG_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  REG_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  REG_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  REG_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  REG_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  REG_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  REG_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  REG_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  REG_9 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  REG_10 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  REG_11 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  REG_12 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  REG_13 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  REG_14 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  REG_15 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  REG_16 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  REG_17 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  REG_18 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  REG_19 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  REG_20 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  REG_21 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  REG_22 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  REG_23 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  REG_24 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  REG_25 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  REG_26 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  REG_27 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  REG_28 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  REG_29 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  REG_30 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  REG_31 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  REG_32 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  REG_33 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  REG_34 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  REG_35 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  REG_36 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  REG_37 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  REG_38 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  REG_39 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  REG_40 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  REG_41 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  REG_42 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  REG_43 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  REG_44 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  REG_45 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  REG_46 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  REG_47 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  REG_48 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  REG_49 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  REG_50 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  REG_51 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  REG_52 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  REG_53 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  REG_54 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  REG_55 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  REG_56 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  REG_57 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  REG_58 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  REG_59 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  REG_60 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  REG_61 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  REG_62 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  REG_63 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  REG_64 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  REG_65 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  REG_66 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  REG_67 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  REG_68 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  REG_69 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  REG_70 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  REG_71 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  REG_72 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  REG_73 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  REG_74 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  REG_75 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  REG_76 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  REG_77 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  REG_78 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  REG_79 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  REG_80 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  REG_81 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  REG_82 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  REG_83 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  REG_84 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  REG_85 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  REG_86 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  REG_87 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  REG_88 = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  REG_89 = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  REG_90 = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  REG_91 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  REG_92 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  REG_93 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  REG_94 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  REG_95 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  REG_96 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  REG_97 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  REG_98 = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  REG_99 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  REG_100 = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  REG_101 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  REG_102 = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  REG_103 = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  REG_104 = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  REG_105 = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  REG_106 = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  REG_107 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  REG_108 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  REG_109 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  REG_110 = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  REG_111 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  REG_112 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  REG_113 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  REG_114 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  REG_115 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  REG_116 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  REG_117 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  REG_118 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  REG_119 = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  REG_120 = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  REG_121 = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  REG_122 = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  REG_123 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  REG_124 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  REG_125 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  REG_126 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  REG_127 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  REG_128 = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  REG_129 = _RAND_129[31:0];
  _RAND_130 = {1{`RANDOM}};
  REG_130 = _RAND_130[31:0];
  _RAND_131 = {1{`RANDOM}};
  REG_131 = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  REG_132 = _RAND_132[31:0];
  _RAND_133 = {1{`RANDOM}};
  REG_133 = _RAND_133[31:0];
  _RAND_134 = {1{`RANDOM}};
  REG_134 = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  REG_135 = _RAND_135[31:0];
  _RAND_136 = {1{`RANDOM}};
  REG_136 = _RAND_136[31:0];
  _RAND_137 = {1{`RANDOM}};
  REG_137 = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  REG_138 = _RAND_138[31:0];
  _RAND_139 = {1{`RANDOM}};
  REG_139 = _RAND_139[31:0];
  _RAND_140 = {1{`RANDOM}};
  REG_140 = _RAND_140[31:0];
  _RAND_141 = {1{`RANDOM}};
  REG_141 = _RAND_141[31:0];
  _RAND_142 = {1{`RANDOM}};
  REG_142 = _RAND_142[31:0];
  _RAND_143 = {1{`RANDOM}};
  REG_143 = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  REG_144 = _RAND_144[31:0];
  _RAND_145 = {1{`RANDOM}};
  REG_145 = _RAND_145[31:0];
  _RAND_146 = {1{`RANDOM}};
  REG_146 = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  REG_147 = _RAND_147[31:0];
  _RAND_148 = {1{`RANDOM}};
  REG_148 = _RAND_148[31:0];
  _RAND_149 = {1{`RANDOM}};
  REG_149 = _RAND_149[31:0];
  _RAND_150 = {1{`RANDOM}};
  REG_150 = _RAND_150[31:0];
  _RAND_151 = {1{`RANDOM}};
  REG_151 = _RAND_151[31:0];
  _RAND_152 = {1{`RANDOM}};
  REG_152 = _RAND_152[31:0];
  _RAND_153 = {1{`RANDOM}};
  REG_153 = _RAND_153[31:0];
  _RAND_154 = {1{`RANDOM}};
  REG_154 = _RAND_154[31:0];
  _RAND_155 = {1{`RANDOM}};
  REG_155 = _RAND_155[31:0];
  _RAND_156 = {1{`RANDOM}};
  REG_156 = _RAND_156[31:0];
  _RAND_157 = {1{`RANDOM}};
  REG_157 = _RAND_157[31:0];
  _RAND_158 = {1{`RANDOM}};
  REG_158 = _RAND_158[31:0];
  _RAND_159 = {1{`RANDOM}};
  REG_159 = _RAND_159[31:0];
  _RAND_160 = {1{`RANDOM}};
  REG_160 = _RAND_160[31:0];
  _RAND_161 = {1{`RANDOM}};
  REG_161 = _RAND_161[31:0];
  _RAND_162 = {1{`RANDOM}};
  REG_162 = _RAND_162[31:0];
  _RAND_163 = {1{`RANDOM}};
  REG_163 = _RAND_163[31:0];
  _RAND_164 = {1{`RANDOM}};
  REG_164 = _RAND_164[31:0];
  _RAND_165 = {1{`RANDOM}};
  REG_165 = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  REG_166 = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  REG_167 = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  REG_168 = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  REG_169 = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  REG_170 = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  REG_171 = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  REG_172 = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  REG_173 = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  REG_174 = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  REG_175 = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  REG_176 = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  REG_177 = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  REG_178 = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  REG_179 = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  REG_180 = _RAND_180[31:0];
  _RAND_181 = {1{`RANDOM}};
  REG_181 = _RAND_181[31:0];
  _RAND_182 = {1{`RANDOM}};
  REG_182 = _RAND_182[31:0];
  _RAND_183 = {1{`RANDOM}};
  REG_183 = _RAND_183[31:0];
  _RAND_184 = {1{`RANDOM}};
  REG_184 = _RAND_184[31:0];
  _RAND_185 = {1{`RANDOM}};
  REG_185 = _RAND_185[31:0];
  _RAND_186 = {1{`RANDOM}};
  REG_186 = _RAND_186[31:0];
  _RAND_187 = {1{`RANDOM}};
  REG_187 = _RAND_187[31:0];
  _RAND_188 = {1{`RANDOM}};
  REG_188 = _RAND_188[31:0];
  _RAND_189 = {1{`RANDOM}};
  REG_189 = _RAND_189[31:0];
  _RAND_190 = {1{`RANDOM}};
  REG_190 = _RAND_190[31:0];
  _RAND_191 = {1{`RANDOM}};
  REG_191 = _RAND_191[31:0];
  _RAND_192 = {1{`RANDOM}};
  REG_192 = _RAND_192[31:0];
  _RAND_193 = {1{`RANDOM}};
  REG_193 = _RAND_193[31:0];
  _RAND_194 = {1{`RANDOM}};
  REG_194 = _RAND_194[31:0];
  _RAND_195 = {1{`RANDOM}};
  REG_195 = _RAND_195[31:0];
  _RAND_196 = {1{`RANDOM}};
  REG_196 = _RAND_196[31:0];
  _RAND_197 = {1{`RANDOM}};
  REG_197 = _RAND_197[31:0];
  _RAND_198 = {1{`RANDOM}};
  REG_198 = _RAND_198[31:0];
  _RAND_199 = {1{`RANDOM}};
  REG_199 = _RAND_199[31:0];
  _RAND_200 = {1{`RANDOM}};
  REG_200 = _RAND_200[31:0];
  _RAND_201 = {1{`RANDOM}};
  REG_201 = _RAND_201[31:0];
  _RAND_202 = {1{`RANDOM}};
  REG_202 = _RAND_202[31:0];
  _RAND_203 = {1{`RANDOM}};
  REG_203 = _RAND_203[31:0];
  _RAND_204 = {1{`RANDOM}};
  REG_204 = _RAND_204[31:0];
  _RAND_205 = {1{`RANDOM}};
  REG_205 = _RAND_205[31:0];
  _RAND_206 = {1{`RANDOM}};
  REG_206 = _RAND_206[31:0];
  _RAND_207 = {1{`RANDOM}};
  REG_207 = _RAND_207[31:0];
  _RAND_208 = {1{`RANDOM}};
  REG_208 = _RAND_208[31:0];
  _RAND_209 = {1{`RANDOM}};
  REG_209 = _RAND_209[31:0];
  _RAND_210 = {1{`RANDOM}};
  REG_210 = _RAND_210[31:0];
  _RAND_211 = {1{`RANDOM}};
  REG_211 = _RAND_211[31:0];
  _RAND_212 = {1{`RANDOM}};
  REG_212 = _RAND_212[31:0];
  _RAND_213 = {1{`RANDOM}};
  REG_213 = _RAND_213[31:0];
  _RAND_214 = {1{`RANDOM}};
  REG_214 = _RAND_214[31:0];
  _RAND_215 = {1{`RANDOM}};
  REG_215 = _RAND_215[31:0];
  _RAND_216 = {1{`RANDOM}};
  REG_216 = _RAND_216[31:0];
  _RAND_217 = {1{`RANDOM}};
  REG_217 = _RAND_217[31:0];
  _RAND_218 = {1{`RANDOM}};
  REG_218 = _RAND_218[31:0];
  _RAND_219 = {1{`RANDOM}};
  REG_219 = _RAND_219[31:0];
  _RAND_220 = {1{`RANDOM}};
  REG_220 = _RAND_220[31:0];
  _RAND_221 = {1{`RANDOM}};
  REG_221 = _RAND_221[31:0];
  _RAND_222 = {1{`RANDOM}};
  REG_222 = _RAND_222[31:0];
  _RAND_223 = {1{`RANDOM}};
  REG_223 = _RAND_223[31:0];
  _RAND_224 = {1{`RANDOM}};
  REG_224 = _RAND_224[31:0];
  _RAND_225 = {1{`RANDOM}};
  REG_225 = _RAND_225[31:0];
  _RAND_226 = {1{`RANDOM}};
  REG_226 = _RAND_226[31:0];
  _RAND_227 = {1{`RANDOM}};
  REG_227 = _RAND_227[31:0];
  _RAND_228 = {1{`RANDOM}};
  REG_228 = _RAND_228[31:0];
  _RAND_229 = {1{`RANDOM}};
  REG_229 = _RAND_229[31:0];
  _RAND_230 = {1{`RANDOM}};
  REG_230 = _RAND_230[31:0];
  _RAND_231 = {1{`RANDOM}};
  REG_231 = _RAND_231[31:0];
  _RAND_232 = {1{`RANDOM}};
  REG_232 = _RAND_232[31:0];
  _RAND_233 = {1{`RANDOM}};
  REG_233 = _RAND_233[31:0];
  _RAND_234 = {1{`RANDOM}};
  REG_234 = _RAND_234[31:0];
  _RAND_235 = {1{`RANDOM}};
  REG_235 = _RAND_235[31:0];
  _RAND_236 = {1{`RANDOM}};
  REG_236 = _RAND_236[31:0];
  _RAND_237 = {1{`RANDOM}};
  REG_237 = _RAND_237[31:0];
  _RAND_238 = {1{`RANDOM}};
  REG_238 = _RAND_238[31:0];
  _RAND_239 = {1{`RANDOM}};
  REG_239 = _RAND_239[31:0];
  _RAND_240 = {1{`RANDOM}};
  REG_240 = _RAND_240[31:0];
  _RAND_241 = {1{`RANDOM}};
  REG_241 = _RAND_241[31:0];
  _RAND_242 = {1{`RANDOM}};
  REG_242 = _RAND_242[31:0];
  _RAND_243 = {1{`RANDOM}};
  REG_243 = _RAND_243[31:0];
  _RAND_244 = {1{`RANDOM}};
  REG_244 = _RAND_244[31:0];
  _RAND_245 = {1{`RANDOM}};
  REG_245 = _RAND_245[31:0];
  _RAND_246 = {1{`RANDOM}};
  REG_246 = _RAND_246[31:0];
  _RAND_247 = {1{`RANDOM}};
  REG_247 = _RAND_247[31:0];
  _RAND_248 = {1{`RANDOM}};
  REG_248 = _RAND_248[31:0];
  _RAND_249 = {1{`RANDOM}};
  REG_249 = _RAND_249[31:0];
  _RAND_250 = {1{`RANDOM}};
  REG_250 = _RAND_250[31:0];
  _RAND_251 = {1{`RANDOM}};
  REG_251 = _RAND_251[31:0];
  _RAND_252 = {1{`RANDOM}};
  REG_252 = _RAND_252[31:0];
  _RAND_253 = {1{`RANDOM}};
  REG_253 = _RAND_253[31:0];
  _RAND_254 = {1{`RANDOM}};
  REG_254 = _RAND_254[31:0];
  _RAND_255 = {1{`RANDOM}};
  REG_255 = _RAND_255[31:0];
  _RAND_256 = {1{`RANDOM}};
  REG_256 = _RAND_256[31:0];
  _RAND_257 = {1{`RANDOM}};
  REG_257 = _RAND_257[31:0];
  _RAND_258 = {1{`RANDOM}};
  REG_258 = _RAND_258[31:0];
  _RAND_259 = {1{`RANDOM}};
  REG_259 = _RAND_259[31:0];
  _RAND_260 = {1{`RANDOM}};
  REG_260 = _RAND_260[31:0];
  _RAND_261 = {1{`RANDOM}};
  REG_261 = _RAND_261[31:0];
  _RAND_262 = {1{`RANDOM}};
  REG_262 = _RAND_262[31:0];
  _RAND_263 = {1{`RANDOM}};
  REG_263 = _RAND_263[31:0];
  _RAND_264 = {1{`RANDOM}};
  REG_264 = _RAND_264[31:0];
  _RAND_265 = {1{`RANDOM}};
  REG_265 = _RAND_265[31:0];
  _RAND_266 = {1{`RANDOM}};
  REG_266 = _RAND_266[31:0];
  _RAND_267 = {1{`RANDOM}};
  REG_267 = _RAND_267[31:0];
  _RAND_268 = {1{`RANDOM}};
  REG_268 = _RAND_268[31:0];
  _RAND_269 = {1{`RANDOM}};
  REG_269 = _RAND_269[31:0];
  _RAND_270 = {1{`RANDOM}};
  REG_270 = _RAND_270[31:0];
  _RAND_271 = {1{`RANDOM}};
  REG_271 = _RAND_271[31:0];
  _RAND_272 = {1{`RANDOM}};
  REG_272 = _RAND_272[31:0];
  _RAND_273 = {1{`RANDOM}};
  REG_273 = _RAND_273[31:0];
  _RAND_274 = {1{`RANDOM}};
  REG_274 = _RAND_274[31:0];
  _RAND_275 = {1{`RANDOM}};
  REG_275 = _RAND_275[31:0];
  _RAND_276 = {1{`RANDOM}};
  REG_276 = _RAND_276[31:0];
  _RAND_277 = {1{`RANDOM}};
  REG_277 = _RAND_277[31:0];
  _RAND_278 = {1{`RANDOM}};
  REG_278 = _RAND_278[31:0];
  _RAND_279 = {1{`RANDOM}};
  REG_279 = _RAND_279[31:0];
  _RAND_280 = {1{`RANDOM}};
  REG_280 = _RAND_280[31:0];
  _RAND_281 = {1{`RANDOM}};
  REG_281 = _RAND_281[31:0];
  _RAND_282 = {1{`RANDOM}};
  REG_282 = _RAND_282[31:0];
  _RAND_283 = {1{`RANDOM}};
  REG_283 = _RAND_283[31:0];
  _RAND_284 = {1{`RANDOM}};
  REG_284 = _RAND_284[31:0];
  _RAND_285 = {1{`RANDOM}};
  REG_285 = _RAND_285[31:0];
  _RAND_286 = {1{`RANDOM}};
  REG_286 = _RAND_286[31:0];
  _RAND_287 = {1{`RANDOM}};
  REG_287 = _RAND_287[31:0];
  _RAND_288 = {1{`RANDOM}};
  REG_288 = _RAND_288[31:0];
  _RAND_289 = {1{`RANDOM}};
  REG_289 = _RAND_289[31:0];
  _RAND_290 = {1{`RANDOM}};
  REG_290 = _RAND_290[31:0];
  _RAND_291 = {1{`RANDOM}};
  REG_291 = _RAND_291[31:0];
  _RAND_292 = {1{`RANDOM}};
  REG_292 = _RAND_292[31:0];
  _RAND_293 = {1{`RANDOM}};
  REG_293 = _RAND_293[31:0];
  _RAND_294 = {1{`RANDOM}};
  REG_294 = _RAND_294[31:0];
  _RAND_295 = {1{`RANDOM}};
  REG_295 = _RAND_295[31:0];
  _RAND_296 = {1{`RANDOM}};
  REG_296 = _RAND_296[31:0];
  _RAND_297 = {1{`RANDOM}};
  REG_297 = _RAND_297[31:0];
  _RAND_298 = {1{`RANDOM}};
  REG_298 = _RAND_298[31:0];
  _RAND_299 = {1{`RANDOM}};
  REG_299 = _RAND_299[31:0];
  _RAND_300 = {1{`RANDOM}};
  REG_300 = _RAND_300[31:0];
  _RAND_301 = {1{`RANDOM}};
  REG_301 = _RAND_301[31:0];
  _RAND_302 = {1{`RANDOM}};
  REG_302 = _RAND_302[31:0];
  _RAND_303 = {1{`RANDOM}};
  REG_303 = _RAND_303[31:0];
  _RAND_304 = {1{`RANDOM}};
  REG_304 = _RAND_304[31:0];
  _RAND_305 = {1{`RANDOM}};
  REG_305 = _RAND_305[31:0];
  _RAND_306 = {1{`RANDOM}};
  REG_306 = _RAND_306[31:0];
  _RAND_307 = {1{`RANDOM}};
  REG_307 = _RAND_307[31:0];
  _RAND_308 = {1{`RANDOM}};
  REG_308 = _RAND_308[31:0];
  _RAND_309 = {1{`RANDOM}};
  REG_309 = _RAND_309[31:0];
  _RAND_310 = {1{`RANDOM}};
  REG_310 = _RAND_310[31:0];
  _RAND_311 = {1{`RANDOM}};
  REG_311 = _RAND_311[31:0];
  _RAND_312 = {1{`RANDOM}};
  REG_312 = _RAND_312[31:0];
  _RAND_313 = {1{`RANDOM}};
  REG_313 = _RAND_313[31:0];
  _RAND_314 = {1{`RANDOM}};
  REG_314 = _RAND_314[31:0];
  _RAND_315 = {1{`RANDOM}};
  REG_315 = _RAND_315[31:0];
  _RAND_316 = {1{`RANDOM}};
  REG_316 = _RAND_316[31:0];
  _RAND_317 = {1{`RANDOM}};
  REG_317 = _RAND_317[31:0];
  _RAND_318 = {1{`RANDOM}};
  REG_318 = _RAND_318[31:0];
  _RAND_319 = {1{`RANDOM}};
  REG_319 = _RAND_319[31:0];
  _RAND_320 = {1{`RANDOM}};
  REG_320 = _RAND_320[31:0];
  _RAND_321 = {1{`RANDOM}};
  REG_321 = _RAND_321[31:0];
  _RAND_322 = {1{`RANDOM}};
  REG_322 = _RAND_322[31:0];
  _RAND_323 = {1{`RANDOM}};
  REG_323 = _RAND_323[31:0];
  _RAND_324 = {1{`RANDOM}};
  REG_324 = _RAND_324[31:0];
  _RAND_325 = {1{`RANDOM}};
  REG_325 = _RAND_325[31:0];
  _RAND_326 = {1{`RANDOM}};
  REG_326 = _RAND_326[31:0];
  _RAND_327 = {1{`RANDOM}};
  REG_327 = _RAND_327[31:0];
  _RAND_328 = {1{`RANDOM}};
  REG_328 = _RAND_328[31:0];
  _RAND_329 = {1{`RANDOM}};
  REG_329 = _RAND_329[31:0];
  _RAND_330 = {1{`RANDOM}};
  REG_330 = _RAND_330[31:0];
  _RAND_331 = {1{`RANDOM}};
  REG_331 = _RAND_331[31:0];
  _RAND_332 = {1{`RANDOM}};
  REG_332 = _RAND_332[31:0];
  _RAND_333 = {1{`RANDOM}};
  REG_333 = _RAND_333[31:0];
  _RAND_334 = {1{`RANDOM}};
  REG_334 = _RAND_334[31:0];
  _RAND_335 = {1{`RANDOM}};
  REG_335 = _RAND_335[31:0];
  _RAND_336 = {1{`RANDOM}};
  REG_336 = _RAND_336[31:0];
  _RAND_337 = {1{`RANDOM}};
  REG_337 = _RAND_337[31:0];
  _RAND_338 = {1{`RANDOM}};
  REG_338 = _RAND_338[31:0];
  _RAND_339 = {1{`RANDOM}};
  REG_339 = _RAND_339[31:0];
  _RAND_340 = {1{`RANDOM}};
  REG_340 = _RAND_340[31:0];
  _RAND_341 = {1{`RANDOM}};
  REG_341 = _RAND_341[31:0];
  _RAND_342 = {1{`RANDOM}};
  REG_342 = _RAND_342[31:0];
  _RAND_343 = {1{`RANDOM}};
  REG_343 = _RAND_343[31:0];
  _RAND_344 = {1{`RANDOM}};
  REG_344 = _RAND_344[31:0];
  _RAND_345 = {1{`RANDOM}};
  REG_345 = _RAND_345[31:0];
  _RAND_346 = {1{`RANDOM}};
  REG_346 = _RAND_346[31:0];
  _RAND_347 = {1{`RANDOM}};
  REG_347 = _RAND_347[31:0];
  _RAND_348 = {1{`RANDOM}};
  REG_348 = _RAND_348[31:0];
  _RAND_349 = {1{`RANDOM}};
  REG_349 = _RAND_349[31:0];
  _RAND_350 = {1{`RANDOM}};
  REG_350 = _RAND_350[31:0];
  _RAND_351 = {1{`RANDOM}};
  REG_351 = _RAND_351[31:0];
  _RAND_352 = {1{`RANDOM}};
  REG_352 = _RAND_352[31:0];
  _RAND_353 = {1{`RANDOM}};
  REG_353 = _RAND_353[31:0];
  _RAND_354 = {1{`RANDOM}};
  REG_354 = _RAND_354[31:0];
  _RAND_355 = {1{`RANDOM}};
  REG_355 = _RAND_355[31:0];
  _RAND_356 = {1{`RANDOM}};
  REG_356 = _RAND_356[31:0];
  _RAND_357 = {1{`RANDOM}};
  REG_357 = _RAND_357[31:0];
  _RAND_358 = {1{`RANDOM}};
  REG_358 = _RAND_358[31:0];
  _RAND_359 = {1{`RANDOM}};
  REG_359 = _RAND_359[31:0];
  _RAND_360 = {1{`RANDOM}};
  REG_360 = _RAND_360[31:0];
  _RAND_361 = {1{`RANDOM}};
  REG_361 = _RAND_361[31:0];
  _RAND_362 = {1{`RANDOM}};
  REG_362 = _RAND_362[31:0];
  _RAND_363 = {1{`RANDOM}};
  REG_363 = _RAND_363[31:0];
  _RAND_364 = {1{`RANDOM}};
  REG_364 = _RAND_364[31:0];
  _RAND_365 = {1{`RANDOM}};
  REG_365 = _RAND_365[31:0];
  _RAND_366 = {1{`RANDOM}};
  REG_366 = _RAND_366[31:0];
  _RAND_367 = {1{`RANDOM}};
  REG_367 = _RAND_367[31:0];
  _RAND_368 = {1{`RANDOM}};
  REG_368 = _RAND_368[31:0];
  _RAND_369 = {1{`RANDOM}};
  REG_369 = _RAND_369[31:0];
  _RAND_370 = {1{`RANDOM}};
  REG_370 = _RAND_370[31:0];
  _RAND_371 = {1{`RANDOM}};
  REG_371 = _RAND_371[31:0];
  _RAND_372 = {1{`RANDOM}};
  REG_372 = _RAND_372[31:0];
  _RAND_373 = {1{`RANDOM}};
  REG_373 = _RAND_373[31:0];
  _RAND_374 = {1{`RANDOM}};
  REG_374 = _RAND_374[31:0];
  _RAND_375 = {1{`RANDOM}};
  REG_375 = _RAND_375[31:0];
  _RAND_376 = {1{`RANDOM}};
  REG_376 = _RAND_376[31:0];
  _RAND_377 = {1{`RANDOM}};
  REG_377 = _RAND_377[31:0];
  _RAND_378 = {1{`RANDOM}};
  REG_378 = _RAND_378[31:0];
  _RAND_379 = {1{`RANDOM}};
  REG_379 = _RAND_379[31:0];
  _RAND_380 = {1{`RANDOM}};
  REG_380 = _RAND_380[31:0];
  _RAND_381 = {1{`RANDOM}};
  REG_381 = _RAND_381[31:0];
  _RAND_382 = {1{`RANDOM}};
  REG_382 = _RAND_382[31:0];
  _RAND_383 = {1{`RANDOM}};
  REG_383 = _RAND_383[31:0];
  _RAND_384 = {1{`RANDOM}};
  REG_384 = _RAND_384[31:0];
  _RAND_385 = {1{`RANDOM}};
  REG_385 = _RAND_385[31:0];
  _RAND_386 = {1{`RANDOM}};
  REG_386 = _RAND_386[31:0];
  _RAND_387 = {1{`RANDOM}};
  REG_387 = _RAND_387[31:0];
  _RAND_388 = {1{`RANDOM}};
  REG_388 = _RAND_388[31:0];
  _RAND_389 = {1{`RANDOM}};
  REG_389 = _RAND_389[31:0];
  _RAND_390 = {1{`RANDOM}};
  REG_390 = _RAND_390[31:0];
  _RAND_391 = {1{`RANDOM}};
  REG_391 = _RAND_391[31:0];
  _RAND_392 = {1{`RANDOM}};
  REG_392 = _RAND_392[31:0];
  _RAND_393 = {1{`RANDOM}};
  REG_393 = _RAND_393[31:0];
  _RAND_394 = {1{`RANDOM}};
  REG_394 = _RAND_394[31:0];
  _RAND_395 = {1{`RANDOM}};
  REG_395 = _RAND_395[31:0];
  _RAND_396 = {1{`RANDOM}};
  REG_396 = _RAND_396[31:0];
  _RAND_397 = {1{`RANDOM}};
  REG_397 = _RAND_397[31:0];
  _RAND_398 = {1{`RANDOM}};
  REG_398 = _RAND_398[31:0];
  _RAND_399 = {1{`RANDOM}};
  REG_399 = _RAND_399[31:0];
  _RAND_400 = {1{`RANDOM}};
  REG_400 = _RAND_400[31:0];
  _RAND_401 = {1{`RANDOM}};
  REG_401 = _RAND_401[31:0];
  _RAND_402 = {1{`RANDOM}};
  REG_402 = _RAND_402[31:0];
  _RAND_403 = {1{`RANDOM}};
  REG_403 = _RAND_403[31:0];
  _RAND_404 = {1{`RANDOM}};
  REG_404 = _RAND_404[31:0];
  _RAND_405 = {1{`RANDOM}};
  REG_405 = _RAND_405[31:0];
  _RAND_406 = {1{`RANDOM}};
  REG_406 = _RAND_406[31:0];
  _RAND_407 = {1{`RANDOM}};
  REG_407 = _RAND_407[31:0];
  _RAND_408 = {1{`RANDOM}};
  REG_408 = _RAND_408[31:0];
  _RAND_409 = {1{`RANDOM}};
  REG_409 = _RAND_409[31:0];
  _RAND_410 = {1{`RANDOM}};
  REG_410 = _RAND_410[31:0];
  _RAND_411 = {1{`RANDOM}};
  REG_411 = _RAND_411[31:0];
  _RAND_412 = {1{`RANDOM}};
  REG_412 = _RAND_412[31:0];
  _RAND_413 = {1{`RANDOM}};
  REG_413 = _RAND_413[31:0];
  _RAND_414 = {1{`RANDOM}};
  REG_414 = _RAND_414[31:0];
  _RAND_415 = {1{`RANDOM}};
  REG_415 = _RAND_415[31:0];
  _RAND_416 = {1{`RANDOM}};
  REG_416 = _RAND_416[31:0];
  _RAND_417 = {1{`RANDOM}};
  REG_417 = _RAND_417[31:0];
  _RAND_418 = {1{`RANDOM}};
  REG_418 = _RAND_418[31:0];
  _RAND_419 = {1{`RANDOM}};
  REG_419 = _RAND_419[31:0];
  _RAND_420 = {1{`RANDOM}};
  REG_420 = _RAND_420[31:0];
  _RAND_421 = {1{`RANDOM}};
  REG_421 = _RAND_421[31:0];
  _RAND_422 = {1{`RANDOM}};
  REG_422 = _RAND_422[31:0];
  _RAND_423 = {1{`RANDOM}};
  REG_423 = _RAND_423[31:0];
  _RAND_424 = {1{`RANDOM}};
  REG_424 = _RAND_424[31:0];
  _RAND_425 = {1{`RANDOM}};
  REG_425 = _RAND_425[31:0];
  _RAND_426 = {1{`RANDOM}};
  REG_426 = _RAND_426[31:0];
  _RAND_427 = {1{`RANDOM}};
  REG_427 = _RAND_427[31:0];
  _RAND_428 = {1{`RANDOM}};
  REG_428 = _RAND_428[31:0];
  _RAND_429 = {1{`RANDOM}};
  REG_429 = _RAND_429[31:0];
  _RAND_430 = {1{`RANDOM}};
  REG_430 = _RAND_430[31:0];
  _RAND_431 = {1{`RANDOM}};
  REG_431 = _RAND_431[31:0];
  _RAND_432 = {1{`RANDOM}};
  REG_432 = _RAND_432[31:0];
  _RAND_433 = {1{`RANDOM}};
  REG_433 = _RAND_433[31:0];
  _RAND_434 = {1{`RANDOM}};
  REG_434 = _RAND_434[31:0];
  _RAND_435 = {1{`RANDOM}};
  REG_435 = _RAND_435[31:0];
  _RAND_436 = {1{`RANDOM}};
  REG_436 = _RAND_436[31:0];
  _RAND_437 = {1{`RANDOM}};
  REG_437 = _RAND_437[31:0];
  _RAND_438 = {1{`RANDOM}};
  REG_438 = _RAND_438[31:0];
  _RAND_439 = {1{`RANDOM}};
  REG_439 = _RAND_439[31:0];
  _RAND_440 = {1{`RANDOM}};
  REG_440 = _RAND_440[31:0];
  _RAND_441 = {1{`RANDOM}};
  REG_441 = _RAND_441[31:0];
  _RAND_442 = {1{`RANDOM}};
  REG_442 = _RAND_442[31:0];
  _RAND_443 = {1{`RANDOM}};
  REG_443 = _RAND_443[31:0];
  _RAND_444 = {1{`RANDOM}};
  REG_444 = _RAND_444[31:0];
  _RAND_445 = {1{`RANDOM}};
  REG_445 = _RAND_445[31:0];
  _RAND_446 = {1{`RANDOM}};
  REG_446 = _RAND_446[31:0];
  _RAND_447 = {1{`RANDOM}};
  REG_447 = _RAND_447[31:0];
  _RAND_448 = {1{`RANDOM}};
  REG_448 = _RAND_448[31:0];
  _RAND_449 = {1{`RANDOM}};
  REG_449 = _RAND_449[31:0];
  _RAND_450 = {1{`RANDOM}};
  REG_450 = _RAND_450[31:0];
  _RAND_451 = {1{`RANDOM}};
  REG_451 = _RAND_451[31:0];
  _RAND_452 = {1{`RANDOM}};
  REG_452 = _RAND_452[31:0];
  _RAND_453 = {1{`RANDOM}};
  REG_453 = _RAND_453[31:0];
  _RAND_454 = {1{`RANDOM}};
  REG_454 = _RAND_454[31:0];
  _RAND_455 = {1{`RANDOM}};
  REG_455 = _RAND_455[31:0];
  _RAND_456 = {1{`RANDOM}};
  REG_456 = _RAND_456[31:0];
  _RAND_457 = {1{`RANDOM}};
  REG_457 = _RAND_457[31:0];
  _RAND_458 = {1{`RANDOM}};
  REG_458 = _RAND_458[31:0];
  _RAND_459 = {1{`RANDOM}};
  REG_459 = _RAND_459[31:0];
  _RAND_460 = {1{`RANDOM}};
  REG_460 = _RAND_460[31:0];
  _RAND_461 = {1{`RANDOM}};
  REG_461 = _RAND_461[31:0];
  _RAND_462 = {1{`RANDOM}};
  REG_462 = _RAND_462[31:0];
  _RAND_463 = {1{`RANDOM}};
  REG_463 = _RAND_463[31:0];
  _RAND_464 = {1{`RANDOM}};
  REG_464 = _RAND_464[31:0];
  _RAND_465 = {1{`RANDOM}};
  REG_465 = _RAND_465[31:0];
  _RAND_466 = {1{`RANDOM}};
  REG_466 = _RAND_466[31:0];
  _RAND_467 = {1{`RANDOM}};
  REG_467 = _RAND_467[31:0];
  _RAND_468 = {1{`RANDOM}};
  REG_468 = _RAND_468[31:0];
  _RAND_469 = {1{`RANDOM}};
  REG_469 = _RAND_469[31:0];
  _RAND_470 = {1{`RANDOM}};
  REG_470 = _RAND_470[31:0];
  _RAND_471 = {1{`RANDOM}};
  REG_471 = _RAND_471[31:0];
  _RAND_472 = {1{`RANDOM}};
  REG_472 = _RAND_472[31:0];
  _RAND_473 = {1{`RANDOM}};
  REG_473 = _RAND_473[31:0];
  _RAND_474 = {1{`RANDOM}};
  REG_474 = _RAND_474[31:0];
  _RAND_475 = {1{`RANDOM}};
  REG_475 = _RAND_475[31:0];
  _RAND_476 = {1{`RANDOM}};
  REG_476 = _RAND_476[31:0];
  _RAND_477 = {1{`RANDOM}};
  REG_477 = _RAND_477[31:0];
  _RAND_478 = {1{`RANDOM}};
  REG_478 = _RAND_478[31:0];
  _RAND_479 = {1{`RANDOM}};
  REG_479 = _RAND_479[31:0];
  _RAND_480 = {1{`RANDOM}};
  REG_480 = _RAND_480[31:0];
  _RAND_481 = {1{`RANDOM}};
  REG_481 = _RAND_481[31:0];
  _RAND_482 = {1{`RANDOM}};
  REG_482 = _RAND_482[31:0];
  _RAND_483 = {1{`RANDOM}};
  REG_483 = _RAND_483[31:0];
  _RAND_484 = {1{`RANDOM}};
  REG_484 = _RAND_484[31:0];
  _RAND_485 = {1{`RANDOM}};
  REG_485 = _RAND_485[31:0];
  _RAND_486 = {1{`RANDOM}};
  REG_486 = _RAND_486[31:0];
  _RAND_487 = {1{`RANDOM}};
  REG_487 = _RAND_487[31:0];
  _RAND_488 = {1{`RANDOM}};
  REG_488 = _RAND_488[31:0];
  _RAND_489 = {1{`RANDOM}};
  REG_489 = _RAND_489[31:0];
  _RAND_490 = {1{`RANDOM}};
  REG_490 = _RAND_490[31:0];
  _RAND_491 = {1{`RANDOM}};
  REG_491 = _RAND_491[31:0];
  _RAND_492 = {1{`RANDOM}};
  REG_492 = _RAND_492[31:0];
  _RAND_493 = {1{`RANDOM}};
  REG_493 = _RAND_493[31:0];
  _RAND_494 = {1{`RANDOM}};
  REG_494 = _RAND_494[31:0];
  _RAND_495 = {1{`RANDOM}};
  REG_495 = _RAND_495[31:0];
  _RAND_496 = {1{`RANDOM}};
  REG_496 = _RAND_496[31:0];
  _RAND_497 = {1{`RANDOM}};
  REG_497 = _RAND_497[31:0];
  _RAND_498 = {1{`RANDOM}};
  REG_498 = _RAND_498[31:0];
  _RAND_499 = {1{`RANDOM}};
  REG_499 = _RAND_499[31:0];
  _RAND_500 = {1{`RANDOM}};
  REG_500 = _RAND_500[31:0];
  _RAND_501 = {1{`RANDOM}};
  REG_501 = _RAND_501[31:0];
  _RAND_502 = {1{`RANDOM}};
  REG_502 = _RAND_502[31:0];
  _RAND_503 = {1{`RANDOM}};
  REG_503 = _RAND_503[31:0];
  _RAND_504 = {1{`RANDOM}};
  REG_504 = _RAND_504[31:0];
  _RAND_505 = {1{`RANDOM}};
  REG_505 = _RAND_505[31:0];
  _RAND_506 = {1{`RANDOM}};
  REG_506 = _RAND_506[31:0];
  _RAND_507 = {1{`RANDOM}};
  REG_507 = _RAND_507[31:0];
  _RAND_508 = {1{`RANDOM}};
  REG_508 = _RAND_508[31:0];
  _RAND_509 = {1{`RANDOM}};
  REG_509 = _RAND_509[31:0];
  _RAND_510 = {1{`RANDOM}};
  REG_510 = _RAND_510[31:0];
  _RAND_511 = {1{`RANDOM}};
  REG_511 = _RAND_511[31:0];
  _RAND_512 = {1{`RANDOM}};
  REG_512 = _RAND_512[31:0];
  _RAND_513 = {1{`RANDOM}};
  REG_513 = _RAND_513[31:0];
  _RAND_514 = {1{`RANDOM}};
  REG_514 = _RAND_514[31:0];
  _RAND_515 = {1{`RANDOM}};
  REG_515 = _RAND_515[31:0];
  _RAND_516 = {1{`RANDOM}};
  REG_516 = _RAND_516[31:0];
  _RAND_517 = {1{`RANDOM}};
  REG_517 = _RAND_517[31:0];
  _RAND_518 = {1{`RANDOM}};
  REG_518 = _RAND_518[31:0];
  _RAND_519 = {1{`RANDOM}};
  REG_519 = _RAND_519[31:0];
  _RAND_520 = {1{`RANDOM}};
  REG_520 = _RAND_520[31:0];
  _RAND_521 = {1{`RANDOM}};
  REG_521 = _RAND_521[31:0];
  _RAND_522 = {1{`RANDOM}};
  REG_522 = _RAND_522[31:0];
  _RAND_523 = {1{`RANDOM}};
  REG_523 = _RAND_523[31:0];
  _RAND_524 = {1{`RANDOM}};
  REG_524 = _RAND_524[31:0];
  _RAND_525 = {1{`RANDOM}};
  REG_525 = _RAND_525[31:0];
  _RAND_526 = {1{`RANDOM}};
  REG_526 = _RAND_526[31:0];
  _RAND_527 = {1{`RANDOM}};
  REG_527 = _RAND_527[31:0];
  _RAND_528 = {1{`RANDOM}};
  REG_528 = _RAND_528[31:0];
  _RAND_529 = {1{`RANDOM}};
  REG_529 = _RAND_529[31:0];
  _RAND_530 = {1{`RANDOM}};
  REG_530 = _RAND_530[31:0];
  _RAND_531 = {1{`RANDOM}};
  REG_531 = _RAND_531[31:0];
  _RAND_532 = {1{`RANDOM}};
  REG_532 = _RAND_532[31:0];
  _RAND_533 = {1{`RANDOM}};
  REG_533 = _RAND_533[31:0];
  _RAND_534 = {1{`RANDOM}};
  REG_534 = _RAND_534[31:0];
  _RAND_535 = {1{`RANDOM}};
  REG_535 = _RAND_535[31:0];
  _RAND_536 = {1{`RANDOM}};
  REG_536 = _RAND_536[31:0];
  _RAND_537 = {1{`RANDOM}};
  REG_537 = _RAND_537[31:0];
  _RAND_538 = {1{`RANDOM}};
  REG_538 = _RAND_538[31:0];
  _RAND_539 = {1{`RANDOM}};
  REG_539 = _RAND_539[31:0];
  _RAND_540 = {1{`RANDOM}};
  REG_540 = _RAND_540[31:0];
  _RAND_541 = {1{`RANDOM}};
  REG_541 = _RAND_541[31:0];
  _RAND_542 = {1{`RANDOM}};
  REG_542 = _RAND_542[31:0];
  _RAND_543 = {1{`RANDOM}};
  REG_543 = _RAND_543[31:0];
  _RAND_544 = {1{`RANDOM}};
  REG_544 = _RAND_544[31:0];
  _RAND_545 = {1{`RANDOM}};
  REG_545 = _RAND_545[31:0];
  _RAND_546 = {1{`RANDOM}};
  REG_546 = _RAND_546[31:0];
  _RAND_547 = {1{`RANDOM}};
  REG_547 = _RAND_547[31:0];
  _RAND_548 = {1{`RANDOM}};
  REG_548 = _RAND_548[31:0];
  _RAND_549 = {1{`RANDOM}};
  REG_549 = _RAND_549[31:0];
  _RAND_550 = {1{`RANDOM}};
  REG_550 = _RAND_550[31:0];
  _RAND_551 = {1{`RANDOM}};
  REG_551 = _RAND_551[31:0];
  _RAND_552 = {1{`RANDOM}};
  REG_552 = _RAND_552[31:0];
  _RAND_553 = {1{`RANDOM}};
  REG_553 = _RAND_553[31:0];
  _RAND_554 = {1{`RANDOM}};
  REG_554 = _RAND_554[31:0];
  _RAND_555 = {1{`RANDOM}};
  REG_555 = _RAND_555[31:0];
  _RAND_556 = {1{`RANDOM}};
  REG_556 = _RAND_556[31:0];
  _RAND_557 = {1{`RANDOM}};
  REG_557 = _RAND_557[31:0];
  _RAND_558 = {1{`RANDOM}};
  REG_558 = _RAND_558[31:0];
  _RAND_559 = {1{`RANDOM}};
  REG_559 = _RAND_559[31:0];
  _RAND_560 = {1{`RANDOM}};
  REG_560 = _RAND_560[31:0];
  _RAND_561 = {1{`RANDOM}};
  REG_561 = _RAND_561[31:0];
  _RAND_562 = {1{`RANDOM}};
  REG_562 = _RAND_562[31:0];
  _RAND_563 = {1{`RANDOM}};
  REG_563 = _RAND_563[31:0];
  _RAND_564 = {1{`RANDOM}};
  REG_564 = _RAND_564[31:0];
  _RAND_565 = {1{`RANDOM}};
  REG_565 = _RAND_565[31:0];
  _RAND_566 = {1{`RANDOM}};
  REG_566 = _RAND_566[31:0];
  _RAND_567 = {1{`RANDOM}};
  REG_567 = _RAND_567[31:0];
  _RAND_568 = {1{`RANDOM}};
  REG_568 = _RAND_568[31:0];
  _RAND_569 = {1{`RANDOM}};
  REG_569 = _RAND_569[31:0];
  _RAND_570 = {1{`RANDOM}};
  REG_570 = _RAND_570[31:0];
  _RAND_571 = {1{`RANDOM}};
  REG_571 = _RAND_571[31:0];
  _RAND_572 = {1{`RANDOM}};
  REG_572 = _RAND_572[31:0];
  _RAND_573 = {1{`RANDOM}};
  REG_573 = _RAND_573[31:0];
  _RAND_574 = {1{`RANDOM}};
  REG_574 = _RAND_574[31:0];
  _RAND_575 = {1{`RANDOM}};
  REG_575 = _RAND_575[31:0];
  _RAND_576 = {1{`RANDOM}};
  REG_576 = _RAND_576[31:0];
  _RAND_577 = {1{`RANDOM}};
  REG_577 = _RAND_577[31:0];
  _RAND_578 = {1{`RANDOM}};
  REG_578 = _RAND_578[31:0];
  _RAND_579 = {1{`RANDOM}};
  REG_579 = _RAND_579[31:0];
  _RAND_580 = {1{`RANDOM}};
  REG_580 = _RAND_580[31:0];
  _RAND_581 = {1{`RANDOM}};
  REG_581 = _RAND_581[31:0];
  _RAND_582 = {1{`RANDOM}};
  REG_582 = _RAND_582[31:0];
  _RAND_583 = {1{`RANDOM}};
  REG_583 = _RAND_583[31:0];
  _RAND_584 = {1{`RANDOM}};
  REG_584 = _RAND_584[31:0];
  _RAND_585 = {1{`RANDOM}};
  REG_585 = _RAND_585[31:0];
  _RAND_586 = {1{`RANDOM}};
  REG_586 = _RAND_586[31:0];
  _RAND_587 = {1{`RANDOM}};
  REG_587 = _RAND_587[31:0];
  _RAND_588 = {1{`RANDOM}};
  REG_588 = _RAND_588[31:0];
  _RAND_589 = {1{`RANDOM}};
  REG_589 = _RAND_589[31:0];
  _RAND_590 = {1{`RANDOM}};
  REG_590 = _RAND_590[31:0];
  _RAND_591 = {1{`RANDOM}};
  REG_591 = _RAND_591[31:0];
  _RAND_592 = {1{`RANDOM}};
  REG_592 = _RAND_592[31:0];
  _RAND_593 = {1{`RANDOM}};
  REG_593 = _RAND_593[31:0];
  _RAND_594 = {1{`RANDOM}};
  REG_594 = _RAND_594[31:0];
  _RAND_595 = {1{`RANDOM}};
  REG_595 = _RAND_595[31:0];
  _RAND_596 = {1{`RANDOM}};
  REG_596 = _RAND_596[31:0];
  _RAND_597 = {1{`RANDOM}};
  REG_597 = _RAND_597[31:0];
  _RAND_598 = {1{`RANDOM}};
  REG_598 = _RAND_598[31:0];
  _RAND_599 = {1{`RANDOM}};
  REG_599 = _RAND_599[31:0];
  _RAND_600 = {1{`RANDOM}};
  REG_600 = _RAND_600[31:0];
  _RAND_601 = {1{`RANDOM}};
  REG_601 = _RAND_601[31:0];
  _RAND_602 = {1{`RANDOM}};
  REG_602 = _RAND_602[31:0];
  _RAND_603 = {1{`RANDOM}};
  REG_603 = _RAND_603[31:0];
  _RAND_604 = {1{`RANDOM}};
  REG_604 = _RAND_604[31:0];
  _RAND_605 = {1{`RANDOM}};
  REG_605 = _RAND_605[31:0];
  _RAND_606 = {1{`RANDOM}};
  REG_606 = _RAND_606[31:0];
  _RAND_607 = {1{`RANDOM}};
  REG_607 = _RAND_607[31:0];
  _RAND_608 = {1{`RANDOM}};
  REG_608 = _RAND_608[31:0];
  _RAND_609 = {1{`RANDOM}};
  REG_609 = _RAND_609[31:0];
  _RAND_610 = {1{`RANDOM}};
  REG_610 = _RAND_610[31:0];
  _RAND_611 = {1{`RANDOM}};
  REG_611 = _RAND_611[31:0];
  _RAND_612 = {1{`RANDOM}};
  REG_612 = _RAND_612[31:0];
  _RAND_613 = {1{`RANDOM}};
  REG_613 = _RAND_613[31:0];
  _RAND_614 = {1{`RANDOM}};
  REG_614 = _RAND_614[31:0];
  _RAND_615 = {1{`RANDOM}};
  REG_615 = _RAND_615[31:0];
  _RAND_616 = {1{`RANDOM}};
  REG_616 = _RAND_616[31:0];
  _RAND_617 = {1{`RANDOM}};
  REG_617 = _RAND_617[31:0];
  _RAND_618 = {1{`RANDOM}};
  REG_618 = _RAND_618[31:0];
  _RAND_619 = {1{`RANDOM}};
  REG_619 = _RAND_619[31:0];
  _RAND_620 = {1{`RANDOM}};
  REG_620 = _RAND_620[31:0];
  _RAND_621 = {1{`RANDOM}};
  REG_621 = _RAND_621[31:0];
  _RAND_622 = {1{`RANDOM}};
  REG_622 = _RAND_622[31:0];
  _RAND_623 = {1{`RANDOM}};
  REG_623 = _RAND_623[31:0];
  _RAND_624 = {1{`RANDOM}};
  REG_624 = _RAND_624[31:0];
  _RAND_625 = {1{`RANDOM}};
  REG_625 = _RAND_625[31:0];
  _RAND_626 = {1{`RANDOM}};
  REG_626 = _RAND_626[31:0];
  _RAND_627 = {1{`RANDOM}};
  REG_627 = _RAND_627[31:0];
  _RAND_628 = {1{`RANDOM}};
  REG_628 = _RAND_628[31:0];
  _RAND_629 = {1{`RANDOM}};
  REG_629 = _RAND_629[31:0];
  _RAND_630 = {1{`RANDOM}};
  REG_630 = _RAND_630[31:0];
  _RAND_631 = {1{`RANDOM}};
  REG_631 = _RAND_631[31:0];
  _RAND_632 = {1{`RANDOM}};
  REG_632 = _RAND_632[31:0];
  _RAND_633 = {1{`RANDOM}};
  REG_633 = _RAND_633[31:0];
  _RAND_634 = {1{`RANDOM}};
  REG_634 = _RAND_634[31:0];
  _RAND_635 = {1{`RANDOM}};
  REG_635 = _RAND_635[31:0];
  _RAND_636 = {1{`RANDOM}};
  REG_636 = _RAND_636[31:0];
  _RAND_637 = {1{`RANDOM}};
  REG_637 = _RAND_637[31:0];
  _RAND_638 = {1{`RANDOM}};
  REG_638 = _RAND_638[31:0];
  _RAND_639 = {1{`RANDOM}};
  REG_639 = _RAND_639[31:0];
  _RAND_640 = {1{`RANDOM}};
  REG_640 = _RAND_640[31:0];
  _RAND_641 = {1{`RANDOM}};
  REG_641 = _RAND_641[31:0];
  _RAND_642 = {1{`RANDOM}};
  REG_642 = _RAND_642[31:0];
  _RAND_643 = {1{`RANDOM}};
  REG_643 = _RAND_643[31:0];
  _RAND_644 = {1{`RANDOM}};
  REG_644 = _RAND_644[31:0];
  _RAND_645 = {1{`RANDOM}};
  REG_645 = _RAND_645[31:0];
  _RAND_646 = {1{`RANDOM}};
  REG_646 = _RAND_646[31:0];
  _RAND_647 = {1{`RANDOM}};
  REG_647 = _RAND_647[31:0];
  _RAND_648 = {1{`RANDOM}};
  REG_648 = _RAND_648[31:0];
  _RAND_649 = {1{`RANDOM}};
  REG_649 = _RAND_649[31:0];
  _RAND_650 = {1{`RANDOM}};
  REG_650 = _RAND_650[31:0];
  _RAND_651 = {1{`RANDOM}};
  REG_651 = _RAND_651[31:0];
  _RAND_652 = {1{`RANDOM}};
  REG_652 = _RAND_652[31:0];
  _RAND_653 = {1{`RANDOM}};
  REG_653 = _RAND_653[31:0];
  _RAND_654 = {1{`RANDOM}};
  REG_654 = _RAND_654[31:0];
  _RAND_655 = {1{`RANDOM}};
  REG_655 = _RAND_655[31:0];
  _RAND_656 = {1{`RANDOM}};
  REG_656 = _RAND_656[31:0];
  _RAND_657 = {1{`RANDOM}};
  REG_657 = _RAND_657[31:0];
  _RAND_658 = {1{`RANDOM}};
  REG_658 = _RAND_658[31:0];
  _RAND_659 = {1{`RANDOM}};
  REG_659 = _RAND_659[31:0];
  _RAND_660 = {1{`RANDOM}};
  REG_660 = _RAND_660[31:0];
  _RAND_661 = {1{`RANDOM}};
  REG_661 = _RAND_661[31:0];
  _RAND_662 = {1{`RANDOM}};
  REG_662 = _RAND_662[31:0];
  _RAND_663 = {1{`RANDOM}};
  REG_663 = _RAND_663[31:0];
  _RAND_664 = {1{`RANDOM}};
  REG_664 = _RAND_664[31:0];
  _RAND_665 = {1{`RANDOM}};
  REG_665 = _RAND_665[31:0];
  _RAND_666 = {1{`RANDOM}};
  REG_666 = _RAND_666[31:0];
  _RAND_667 = {1{`RANDOM}};
  REG_667 = _RAND_667[31:0];
  _RAND_668 = {1{`RANDOM}};
  REG_668 = _RAND_668[31:0];
  _RAND_669 = {1{`RANDOM}};
  REG_669 = _RAND_669[31:0];
  _RAND_670 = {1{`RANDOM}};
  REG_670 = _RAND_670[31:0];
  _RAND_671 = {1{`RANDOM}};
  REG_671 = _RAND_671[31:0];
  _RAND_672 = {1{`RANDOM}};
  REG_672 = _RAND_672[31:0];
  _RAND_673 = {1{`RANDOM}};
  REG_673 = _RAND_673[31:0];
  _RAND_674 = {1{`RANDOM}};
  REG_674 = _RAND_674[31:0];
  _RAND_675 = {1{`RANDOM}};
  REG_675 = _RAND_675[31:0];
  _RAND_676 = {1{`RANDOM}};
  REG_676 = _RAND_676[31:0];
  _RAND_677 = {1{`RANDOM}};
  REG_677 = _RAND_677[31:0];
  _RAND_678 = {1{`RANDOM}};
  REG_678 = _RAND_678[31:0];
  _RAND_679 = {1{`RANDOM}};
  REG_679 = _RAND_679[31:0];
  _RAND_680 = {1{`RANDOM}};
  REG_680 = _RAND_680[31:0];
  _RAND_681 = {1{`RANDOM}};
  REG_681 = _RAND_681[31:0];
  _RAND_682 = {1{`RANDOM}};
  REG_682 = _RAND_682[31:0];
  _RAND_683 = {1{`RANDOM}};
  REG_683 = _RAND_683[31:0];
  _RAND_684 = {1{`RANDOM}};
  REG_684 = _RAND_684[31:0];
  _RAND_685 = {1{`RANDOM}};
  REG_685 = _RAND_685[31:0];
  _RAND_686 = {1{`RANDOM}};
  REG_686 = _RAND_686[31:0];
  _RAND_687 = {1{`RANDOM}};
  REG_687 = _RAND_687[31:0];
  _RAND_688 = {1{`RANDOM}};
  REG_688 = _RAND_688[31:0];
  _RAND_689 = {1{`RANDOM}};
  REG_689 = _RAND_689[31:0];
  _RAND_690 = {1{`RANDOM}};
  REG_690 = _RAND_690[31:0];
  _RAND_691 = {1{`RANDOM}};
  REG_691 = _RAND_691[31:0];
  _RAND_692 = {1{`RANDOM}};
  REG_692 = _RAND_692[31:0];
  _RAND_693 = {1{`RANDOM}};
  REG_693 = _RAND_693[31:0];
  _RAND_694 = {1{`RANDOM}};
  REG_694 = _RAND_694[31:0];
  _RAND_695 = {1{`RANDOM}};
  REG_695 = _RAND_695[31:0];
  _RAND_696 = {1{`RANDOM}};
  REG_696 = _RAND_696[31:0];
  _RAND_697 = {1{`RANDOM}};
  REG_697 = _RAND_697[31:0];
  _RAND_698 = {1{`RANDOM}};
  REG_698 = _RAND_698[31:0];
  _RAND_699 = {1{`RANDOM}};
  REG_699 = _RAND_699[31:0];
  _RAND_700 = {1{`RANDOM}};
  REG_700 = _RAND_700[31:0];
  _RAND_701 = {1{`RANDOM}};
  REG_701 = _RAND_701[31:0];
  _RAND_702 = {1{`RANDOM}};
  REG_702 = _RAND_702[31:0];
  _RAND_703 = {1{`RANDOM}};
  REG_703 = _RAND_703[31:0];
  _RAND_704 = {1{`RANDOM}};
  REG_704 = _RAND_704[31:0];
  _RAND_705 = {1{`RANDOM}};
  REG_705 = _RAND_705[31:0];
  _RAND_706 = {1{`RANDOM}};
  REG_706 = _RAND_706[31:0];
  _RAND_707 = {1{`RANDOM}};
  REG_707 = _RAND_707[31:0];
  _RAND_708 = {1{`RANDOM}};
  REG_708 = _RAND_708[31:0];
  _RAND_709 = {1{`RANDOM}};
  REG_709 = _RAND_709[31:0];
  _RAND_710 = {1{`RANDOM}};
  REG_710 = _RAND_710[31:0];
  _RAND_711 = {1{`RANDOM}};
  REG_711 = _RAND_711[31:0];
  _RAND_712 = {1{`RANDOM}};
  REG_712 = _RAND_712[31:0];
  _RAND_713 = {1{`RANDOM}};
  REG_713 = _RAND_713[31:0];
  _RAND_714 = {1{`RANDOM}};
  REG_714 = _RAND_714[31:0];
  _RAND_715 = {1{`RANDOM}};
  REG_715 = _RAND_715[31:0];
  _RAND_716 = {1{`RANDOM}};
  REG_716 = _RAND_716[31:0];
  _RAND_717 = {1{`RANDOM}};
  REG_717 = _RAND_717[31:0];
  _RAND_718 = {1{`RANDOM}};
  REG_718 = _RAND_718[31:0];
  _RAND_719 = {1{`RANDOM}};
  REG_719 = _RAND_719[31:0];
  _RAND_720 = {1{`RANDOM}};
  REG_720 = _RAND_720[31:0];
  _RAND_721 = {1{`RANDOM}};
  REG_721 = _RAND_721[31:0];
  _RAND_722 = {1{`RANDOM}};
  REG_722 = _RAND_722[31:0];
  _RAND_723 = {1{`RANDOM}};
  REG_723 = _RAND_723[31:0];
  _RAND_724 = {1{`RANDOM}};
  REG_724 = _RAND_724[31:0];
  _RAND_725 = {1{`RANDOM}};
  REG_725 = _RAND_725[31:0];
  _RAND_726 = {1{`RANDOM}};
  REG_726 = _RAND_726[31:0];
  _RAND_727 = {1{`RANDOM}};
  REG_727 = _RAND_727[31:0];
  _RAND_728 = {1{`RANDOM}};
  REG_728 = _RAND_728[31:0];
  _RAND_729 = {1{`RANDOM}};
  REG_729 = _RAND_729[31:0];
  _RAND_730 = {1{`RANDOM}};
  REG_730 = _RAND_730[31:0];
  _RAND_731 = {1{`RANDOM}};
  REG_731 = _RAND_731[31:0];
  _RAND_732 = {1{`RANDOM}};
  REG_732 = _RAND_732[31:0];
  _RAND_733 = {1{`RANDOM}};
  REG_733 = _RAND_733[31:0];
  _RAND_734 = {1{`RANDOM}};
  REG_734 = _RAND_734[31:0];
  _RAND_735 = {1{`RANDOM}};
  REG_735 = _RAND_735[31:0];
  _RAND_736 = {1{`RANDOM}};
  REG_736 = _RAND_736[31:0];
  _RAND_737 = {1{`RANDOM}};
  REG_737 = _RAND_737[31:0];
  _RAND_738 = {1{`RANDOM}};
  REG_738 = _RAND_738[31:0];
  _RAND_739 = {1{`RANDOM}};
  REG_739 = _RAND_739[31:0];
  _RAND_740 = {1{`RANDOM}};
  REG_740 = _RAND_740[31:0];
  _RAND_741 = {1{`RANDOM}};
  REG_741 = _RAND_741[31:0];
  _RAND_742 = {1{`RANDOM}};
  REG_742 = _RAND_742[31:0];
  _RAND_743 = {1{`RANDOM}};
  REG_743 = _RAND_743[31:0];
  _RAND_744 = {1{`RANDOM}};
  REG_744 = _RAND_744[31:0];
  _RAND_745 = {1{`RANDOM}};
  REG_745 = _RAND_745[31:0];
  _RAND_746 = {1{`RANDOM}};
  REG_746 = _RAND_746[31:0];
  _RAND_747 = {1{`RANDOM}};
  REG_747 = _RAND_747[31:0];
  _RAND_748 = {1{`RANDOM}};
  REG_748 = _RAND_748[31:0];
  _RAND_749 = {1{`RANDOM}};
  REG_749 = _RAND_749[31:0];
  _RAND_750 = {1{`RANDOM}};
  REG_750 = _RAND_750[31:0];
  _RAND_751 = {1{`RANDOM}};
  REG_751 = _RAND_751[31:0];
  _RAND_752 = {1{`RANDOM}};
  REG_752 = _RAND_752[31:0];
  _RAND_753 = {1{`RANDOM}};
  REG_753 = _RAND_753[31:0];
  _RAND_754 = {1{`RANDOM}};
  REG_754 = _RAND_754[31:0];
  _RAND_755 = {1{`RANDOM}};
  REG_755 = _RAND_755[31:0];
  _RAND_756 = {1{`RANDOM}};
  REG_756 = _RAND_756[31:0];
  _RAND_757 = {1{`RANDOM}};
  REG_757 = _RAND_757[31:0];
  _RAND_758 = {1{`RANDOM}};
  REG_758 = _RAND_758[31:0];
  _RAND_759 = {1{`RANDOM}};
  REG_759 = _RAND_759[31:0];
  _RAND_760 = {1{`RANDOM}};
  REG_760 = _RAND_760[31:0];
  _RAND_761 = {1{`RANDOM}};
  REG_761 = _RAND_761[31:0];
  _RAND_762 = {1{`RANDOM}};
  REG_762 = _RAND_762[31:0];
  _RAND_763 = {1{`RANDOM}};
  REG_763 = _RAND_763[31:0];
  _RAND_764 = {1{`RANDOM}};
  REG_764 = _RAND_764[31:0];
  _RAND_765 = {1{`RANDOM}};
  REG_765 = _RAND_765[31:0];
  _RAND_766 = {1{`RANDOM}};
  REG_766 = _RAND_766[31:0];
  _RAND_767 = {1{`RANDOM}};
  REG_767 = _RAND_767[31:0];
  _RAND_768 = {1{`RANDOM}};
  REG_768 = _RAND_768[31:0];
  _RAND_769 = {1{`RANDOM}};
  REG_769 = _RAND_769[31:0];
  _RAND_770 = {1{`RANDOM}};
  REG_770 = _RAND_770[31:0];
  _RAND_771 = {1{`RANDOM}};
  REG_771 = _RAND_771[31:0];
  _RAND_772 = {1{`RANDOM}};
  REG_772 = _RAND_772[31:0];
  _RAND_773 = {1{`RANDOM}};
  REG_773 = _RAND_773[31:0];
  _RAND_774 = {1{`RANDOM}};
  REG_774 = _RAND_774[31:0];
  _RAND_775 = {1{`RANDOM}};
  REG_775 = _RAND_775[31:0];
  _RAND_776 = {1{`RANDOM}};
  REG_776 = _RAND_776[31:0];
  _RAND_777 = {1{`RANDOM}};
  REG_777 = _RAND_777[31:0];
  _RAND_778 = {1{`RANDOM}};
  REG_778 = _RAND_778[31:0];
  _RAND_779 = {1{`RANDOM}};
  REG_779 = _RAND_779[31:0];
  _RAND_780 = {1{`RANDOM}};
  REG_780 = _RAND_780[31:0];
  _RAND_781 = {1{`RANDOM}};
  REG_781 = _RAND_781[31:0];
  _RAND_782 = {1{`RANDOM}};
  REG_782 = _RAND_782[31:0];
  _RAND_783 = {1{`RANDOM}};
  REG_783 = _RAND_783[31:0];
  _RAND_784 = {1{`RANDOM}};
  REG_784 = _RAND_784[31:0];
  _RAND_785 = {1{`RANDOM}};
  REG_785 = _RAND_785[31:0];
  _RAND_786 = {1{`RANDOM}};
  REG_786 = _RAND_786[31:0];
  _RAND_787 = {1{`RANDOM}};
  REG_787 = _RAND_787[31:0];
  _RAND_788 = {1{`RANDOM}};
  REG_788 = _RAND_788[31:0];
  _RAND_789 = {1{`RANDOM}};
  REG_789 = _RAND_789[31:0];
  _RAND_790 = {1{`RANDOM}};
  REG_790 = _RAND_790[31:0];
  _RAND_791 = {1{`RANDOM}};
  REG_791 = _RAND_791[31:0];
  _RAND_792 = {1{`RANDOM}};
  REG_792 = _RAND_792[31:0];
  _RAND_793 = {1{`RANDOM}};
  REG_793 = _RAND_793[31:0];
  _RAND_794 = {1{`RANDOM}};
  REG_794 = _RAND_794[31:0];
  _RAND_795 = {1{`RANDOM}};
  REG_795 = _RAND_795[31:0];
  _RAND_796 = {1{`RANDOM}};
  REG_796 = _RAND_796[31:0];
  _RAND_797 = {1{`RANDOM}};
  REG_797 = _RAND_797[31:0];
  _RAND_798 = {1{`RANDOM}};
  REG_798 = _RAND_798[31:0];
  _RAND_799 = {1{`RANDOM}};
  REG_799 = _RAND_799[31:0];
  _RAND_800 = {1{`RANDOM}};
  REG_800 = _RAND_800[31:0];
  _RAND_801 = {1{`RANDOM}};
  REG_801 = _RAND_801[31:0];
  _RAND_802 = {1{`RANDOM}};
  REG_802 = _RAND_802[31:0];
  _RAND_803 = {1{`RANDOM}};
  REG_803 = _RAND_803[31:0];
  _RAND_804 = {1{`RANDOM}};
  REG_804 = _RAND_804[31:0];
  _RAND_805 = {1{`RANDOM}};
  REG_805 = _RAND_805[31:0];
  _RAND_806 = {1{`RANDOM}};
  REG_806 = _RAND_806[31:0];
  _RAND_807 = {1{`RANDOM}};
  REG_807 = _RAND_807[31:0];
  _RAND_808 = {1{`RANDOM}};
  REG_808 = _RAND_808[31:0];
  _RAND_809 = {1{`RANDOM}};
  REG_809 = _RAND_809[31:0];
  _RAND_810 = {1{`RANDOM}};
  REG_810 = _RAND_810[31:0];
  _RAND_811 = {1{`RANDOM}};
  REG_811 = _RAND_811[31:0];
  _RAND_812 = {1{`RANDOM}};
  REG_812 = _RAND_812[31:0];
  _RAND_813 = {1{`RANDOM}};
  REG_813 = _RAND_813[31:0];
  _RAND_814 = {1{`RANDOM}};
  REG_814 = _RAND_814[31:0];
  _RAND_815 = {1{`RANDOM}};
  REG_815 = _RAND_815[31:0];
  _RAND_816 = {1{`RANDOM}};
  REG_816 = _RAND_816[31:0];
  _RAND_817 = {1{`RANDOM}};
  REG_817 = _RAND_817[31:0];
  _RAND_818 = {1{`RANDOM}};
  REG_818 = _RAND_818[31:0];
  _RAND_819 = {1{`RANDOM}};
  REG_819 = _RAND_819[31:0];
  _RAND_820 = {1{`RANDOM}};
  REG_820 = _RAND_820[31:0];
  _RAND_821 = {1{`RANDOM}};
  REG_821 = _RAND_821[31:0];
  _RAND_822 = {1{`RANDOM}};
  REG_822 = _RAND_822[31:0];
  _RAND_823 = {1{`RANDOM}};
  REG_823 = _RAND_823[31:0];
  _RAND_824 = {1{`RANDOM}};
  REG_824 = _RAND_824[31:0];
  _RAND_825 = {1{`RANDOM}};
  REG_825 = _RAND_825[31:0];
  _RAND_826 = {1{`RANDOM}};
  REG_826 = _RAND_826[31:0];
  _RAND_827 = {1{`RANDOM}};
  REG_827 = _RAND_827[31:0];
  _RAND_828 = {1{`RANDOM}};
  REG_828 = _RAND_828[31:0];
  _RAND_829 = {1{`RANDOM}};
  REG_829 = _RAND_829[31:0];
  _RAND_830 = {1{`RANDOM}};
  REG_830 = _RAND_830[31:0];
  _RAND_831 = {1{`RANDOM}};
  REG_831 = _RAND_831[31:0];
  _RAND_832 = {1{`RANDOM}};
  REG_832 = _RAND_832[31:0];
  _RAND_833 = {1{`RANDOM}};
  REG_833 = _RAND_833[31:0];
  _RAND_834 = {1{`RANDOM}};
  REG_834 = _RAND_834[31:0];
  _RAND_835 = {1{`RANDOM}};
  REG_835 = _RAND_835[31:0];
  _RAND_836 = {1{`RANDOM}};
  REG_836 = _RAND_836[31:0];
  _RAND_837 = {1{`RANDOM}};
  REG_837 = _RAND_837[31:0];
  _RAND_838 = {1{`RANDOM}};
  REG_838 = _RAND_838[31:0];
  _RAND_839 = {1{`RANDOM}};
  REG_839 = _RAND_839[31:0];
  _RAND_840 = {1{`RANDOM}};
  REG_840 = _RAND_840[31:0];
  _RAND_841 = {1{`RANDOM}};
  REG_841 = _RAND_841[31:0];
  _RAND_842 = {1{`RANDOM}};
  REG_842 = _RAND_842[31:0];
  _RAND_843 = {1{`RANDOM}};
  REG_843 = _RAND_843[31:0];
  _RAND_844 = {1{`RANDOM}};
  REG_844 = _RAND_844[31:0];
  _RAND_845 = {1{`RANDOM}};
  REG_845 = _RAND_845[31:0];
  _RAND_846 = {1{`RANDOM}};
  REG_846 = _RAND_846[31:0];
  _RAND_847 = {1{`RANDOM}};
  REG_847 = _RAND_847[31:0];
  _RAND_848 = {1{`RANDOM}};
  REG_848 = _RAND_848[31:0];
  _RAND_849 = {1{`RANDOM}};
  REG_849 = _RAND_849[31:0];
  _RAND_850 = {1{`RANDOM}};
  REG_850 = _RAND_850[31:0];
  _RAND_851 = {1{`RANDOM}};
  REG_851 = _RAND_851[31:0];
  _RAND_852 = {1{`RANDOM}};
  REG_852 = _RAND_852[31:0];
  _RAND_853 = {1{`RANDOM}};
  REG_853 = _RAND_853[31:0];
  _RAND_854 = {1{`RANDOM}};
  REG_854 = _RAND_854[31:0];
  _RAND_855 = {1{`RANDOM}};
  REG_855 = _RAND_855[31:0];
  _RAND_856 = {1{`RANDOM}};
  REG_856 = _RAND_856[31:0];
  _RAND_857 = {1{`RANDOM}};
  REG_857 = _RAND_857[31:0];
  _RAND_858 = {1{`RANDOM}};
  REG_858 = _RAND_858[31:0];
  _RAND_859 = {1{`RANDOM}};
  REG_859 = _RAND_859[31:0];
  _RAND_860 = {1{`RANDOM}};
  REG_860 = _RAND_860[31:0];
  _RAND_861 = {1{`RANDOM}};
  REG_861 = _RAND_861[31:0];
  _RAND_862 = {1{`RANDOM}};
  REG_862 = _RAND_862[31:0];
  _RAND_863 = {1{`RANDOM}};
  REG_863 = _RAND_863[31:0];
  _RAND_864 = {1{`RANDOM}};
  REG_864 = _RAND_864[31:0];
  _RAND_865 = {1{`RANDOM}};
  REG_865 = _RAND_865[31:0];
  _RAND_866 = {1{`RANDOM}};
  REG_866 = _RAND_866[31:0];
  _RAND_867 = {1{`RANDOM}};
  REG_867 = _RAND_867[31:0];
  _RAND_868 = {1{`RANDOM}};
  REG_868 = _RAND_868[31:0];
  _RAND_869 = {1{`RANDOM}};
  REG_869 = _RAND_869[31:0];
  _RAND_870 = {1{`RANDOM}};
  REG_870 = _RAND_870[31:0];
  _RAND_871 = {1{`RANDOM}};
  REG_871 = _RAND_871[31:0];
  _RAND_872 = {1{`RANDOM}};
  REG_872 = _RAND_872[31:0];
  _RAND_873 = {1{`RANDOM}};
  REG_873 = _RAND_873[31:0];
  _RAND_874 = {1{`RANDOM}};
  REG_874 = _RAND_874[31:0];
  _RAND_875 = {1{`RANDOM}};
  REG_875 = _RAND_875[31:0];
  _RAND_876 = {1{`RANDOM}};
  REG_876 = _RAND_876[31:0];
  _RAND_877 = {1{`RANDOM}};
  REG_877 = _RAND_877[31:0];
  _RAND_878 = {1{`RANDOM}};
  REG_878 = _RAND_878[31:0];
  _RAND_879 = {1{`RANDOM}};
  REG_879 = _RAND_879[31:0];
  _RAND_880 = {1{`RANDOM}};
  REG_880 = _RAND_880[31:0];
  _RAND_881 = {1{`RANDOM}};
  REG_881 = _RAND_881[31:0];
  _RAND_882 = {1{`RANDOM}};
  REG_882 = _RAND_882[31:0];
  _RAND_883 = {1{`RANDOM}};
  REG_883 = _RAND_883[31:0];
  _RAND_884 = {1{`RANDOM}};
  REG_884 = _RAND_884[31:0];
  _RAND_885 = {1{`RANDOM}};
  REG_885 = _RAND_885[31:0];
  _RAND_886 = {1{`RANDOM}};
  REG_886 = _RAND_886[31:0];
  _RAND_887 = {1{`RANDOM}};
  REG_887 = _RAND_887[31:0];
  _RAND_888 = {1{`RANDOM}};
  REG_888 = _RAND_888[31:0];
  _RAND_889 = {1{`RANDOM}};
  REG_889 = _RAND_889[31:0];
  _RAND_890 = {1{`RANDOM}};
  REG_890 = _RAND_890[31:0];
  _RAND_891 = {1{`RANDOM}};
  REG_891 = _RAND_891[31:0];
  _RAND_892 = {1{`RANDOM}};
  REG_892 = _RAND_892[31:0];
  _RAND_893 = {1{`RANDOM}};
  REG_893 = _RAND_893[31:0];
  _RAND_894 = {1{`RANDOM}};
  REG_894 = _RAND_894[31:0];
  _RAND_895 = {1{`RANDOM}};
  REG_895 = _RAND_895[31:0];
  _RAND_896 = {1{`RANDOM}};
  REG_896 = _RAND_896[31:0];
  _RAND_897 = {1{`RANDOM}};
  REG_897 = _RAND_897[31:0];
  _RAND_898 = {1{`RANDOM}};
  REG_898 = _RAND_898[31:0];
  _RAND_899 = {1{`RANDOM}};
  REG_899 = _RAND_899[31:0];
  _RAND_900 = {1{`RANDOM}};
  REG_900 = _RAND_900[31:0];
  _RAND_901 = {1{`RANDOM}};
  REG_901 = _RAND_901[31:0];
  _RAND_902 = {1{`RANDOM}};
  REG_902 = _RAND_902[31:0];
  _RAND_903 = {1{`RANDOM}};
  REG_903 = _RAND_903[31:0];
  _RAND_904 = {1{`RANDOM}};
  REG_904 = _RAND_904[31:0];
  _RAND_905 = {1{`RANDOM}};
  REG_905 = _RAND_905[31:0];
  _RAND_906 = {1{`RANDOM}};
  REG_906 = _RAND_906[31:0];
  _RAND_907 = {1{`RANDOM}};
  REG_907 = _RAND_907[31:0];
  _RAND_908 = {1{`RANDOM}};
  REG_908 = _RAND_908[31:0];
  _RAND_909 = {1{`RANDOM}};
  REG_909 = _RAND_909[31:0];
  _RAND_910 = {1{`RANDOM}};
  REG_910 = _RAND_910[31:0];
  _RAND_911 = {1{`RANDOM}};
  REG_911 = _RAND_911[31:0];
  _RAND_912 = {1{`RANDOM}};
  REG_912 = _RAND_912[31:0];
  _RAND_913 = {1{`RANDOM}};
  REG_913 = _RAND_913[31:0];
  _RAND_914 = {1{`RANDOM}};
  REG_914 = _RAND_914[31:0];
  _RAND_915 = {1{`RANDOM}};
  REG_915 = _RAND_915[31:0];
  _RAND_916 = {1{`RANDOM}};
  REG_916 = _RAND_916[31:0];
  _RAND_917 = {1{`RANDOM}};
  REG_917 = _RAND_917[31:0];
  _RAND_918 = {1{`RANDOM}};
  REG_918 = _RAND_918[31:0];
  _RAND_919 = {1{`RANDOM}};
  REG_919 = _RAND_919[31:0];
  _RAND_920 = {1{`RANDOM}};
  REG_920 = _RAND_920[31:0];
  _RAND_921 = {1{`RANDOM}};
  REG_921 = _RAND_921[31:0];
  _RAND_922 = {1{`RANDOM}};
  REG_922 = _RAND_922[31:0];
  _RAND_923 = {1{`RANDOM}};
  REG_923 = _RAND_923[31:0];
  _RAND_924 = {1{`RANDOM}};
  REG_924 = _RAND_924[31:0];
  _RAND_925 = {1{`RANDOM}};
  REG_925 = _RAND_925[31:0];
  _RAND_926 = {1{`RANDOM}};
  REG_926 = _RAND_926[31:0];
  _RAND_927 = {1{`RANDOM}};
  REG_927 = _RAND_927[31:0];
  _RAND_928 = {1{`RANDOM}};
  REG_928 = _RAND_928[31:0];
  _RAND_929 = {1{`RANDOM}};
  REG_929 = _RAND_929[31:0];
  _RAND_930 = {1{`RANDOM}};
  REG_930 = _RAND_930[31:0];
  _RAND_931 = {1{`RANDOM}};
  REG_931 = _RAND_931[31:0];
  _RAND_932 = {1{`RANDOM}};
  REG_932 = _RAND_932[31:0];
  _RAND_933 = {1{`RANDOM}};
  REG_933 = _RAND_933[31:0];
  _RAND_934 = {1{`RANDOM}};
  REG_934 = _RAND_934[31:0];
  _RAND_935 = {1{`RANDOM}};
  REG_935 = _RAND_935[31:0];
  _RAND_936 = {1{`RANDOM}};
  REG_936 = _RAND_936[31:0];
  _RAND_937 = {1{`RANDOM}};
  REG_937 = _RAND_937[31:0];
  _RAND_938 = {1{`RANDOM}};
  REG_938 = _RAND_938[31:0];
  _RAND_939 = {1{`RANDOM}};
  REG_939 = _RAND_939[31:0];
  _RAND_940 = {1{`RANDOM}};
  REG_940 = _RAND_940[31:0];
  _RAND_941 = {1{`RANDOM}};
  REG_941 = _RAND_941[31:0];
  _RAND_942 = {1{`RANDOM}};
  REG_942 = _RAND_942[31:0];
  _RAND_943 = {1{`RANDOM}};
  REG_943 = _RAND_943[31:0];
  _RAND_944 = {1{`RANDOM}};
  REG_944 = _RAND_944[31:0];
  _RAND_945 = {1{`RANDOM}};
  REG_945 = _RAND_945[31:0];
  _RAND_946 = {1{`RANDOM}};
  REG_946 = _RAND_946[31:0];
  _RAND_947 = {1{`RANDOM}};
  REG_947 = _RAND_947[31:0];
  _RAND_948 = {1{`RANDOM}};
  REG_948 = _RAND_948[31:0];
  _RAND_949 = {1{`RANDOM}};
  REG_949 = _RAND_949[31:0];
  _RAND_950 = {1{`RANDOM}};
  REG_950 = _RAND_950[31:0];
  _RAND_951 = {1{`RANDOM}};
  REG_951 = _RAND_951[31:0];
  _RAND_952 = {1{`RANDOM}};
  REG_952 = _RAND_952[31:0];
  _RAND_953 = {1{`RANDOM}};
  REG_953 = _RAND_953[31:0];
  _RAND_954 = {1{`RANDOM}};
  REG_954 = _RAND_954[31:0];
  _RAND_955 = {1{`RANDOM}};
  REG_955 = _RAND_955[31:0];
  _RAND_956 = {1{`RANDOM}};
  REG_956 = _RAND_956[31:0];
  _RAND_957 = {1{`RANDOM}};
  REG_957 = _RAND_957[31:0];
  _RAND_958 = {1{`RANDOM}};
  REG_958 = _RAND_958[31:0];
  _RAND_959 = {1{`RANDOM}};
  REG_959 = _RAND_959[31:0];
  _RAND_960 = {1{`RANDOM}};
  REG_960 = _RAND_960[31:0];
  _RAND_961 = {1{`RANDOM}};
  REG_961 = _RAND_961[31:0];
  _RAND_962 = {1{`RANDOM}};
  REG_962 = _RAND_962[31:0];
  _RAND_963 = {1{`RANDOM}};
  REG_963 = _RAND_963[31:0];
  _RAND_964 = {1{`RANDOM}};
  REG_964 = _RAND_964[31:0];
  _RAND_965 = {1{`RANDOM}};
  REG_965 = _RAND_965[31:0];
  _RAND_966 = {1{`RANDOM}};
  REG_966 = _RAND_966[31:0];
  _RAND_967 = {1{`RANDOM}};
  REG_967 = _RAND_967[31:0];
  _RAND_968 = {1{`RANDOM}};
  REG_968 = _RAND_968[31:0];
  _RAND_969 = {1{`RANDOM}};
  REG_969 = _RAND_969[31:0];
  _RAND_970 = {1{`RANDOM}};
  REG_970 = _RAND_970[31:0];
  _RAND_971 = {1{`RANDOM}};
  REG_971 = _RAND_971[31:0];
  _RAND_972 = {1{`RANDOM}};
  REG_972 = _RAND_972[31:0];
  _RAND_973 = {1{`RANDOM}};
  REG_973 = _RAND_973[31:0];
  _RAND_974 = {1{`RANDOM}};
  REG_974 = _RAND_974[31:0];
  _RAND_975 = {1{`RANDOM}};
  REG_975 = _RAND_975[31:0];
  _RAND_976 = {1{`RANDOM}};
  REG_976 = _RAND_976[31:0];
  _RAND_977 = {1{`RANDOM}};
  REG_977 = _RAND_977[31:0];
  _RAND_978 = {1{`RANDOM}};
  REG_978 = _RAND_978[31:0];
  _RAND_979 = {1{`RANDOM}};
  REG_979 = _RAND_979[31:0];
  _RAND_980 = {1{`RANDOM}};
  REG_980 = _RAND_980[31:0];
  _RAND_981 = {1{`RANDOM}};
  REG_981 = _RAND_981[31:0];
  _RAND_982 = {1{`RANDOM}};
  REG_982 = _RAND_982[31:0];
  _RAND_983 = {1{`RANDOM}};
  REG_983 = _RAND_983[31:0];
  _RAND_984 = {1{`RANDOM}};
  REG_984 = _RAND_984[31:0];
  _RAND_985 = {1{`RANDOM}};
  REG_985 = _RAND_985[31:0];
  _RAND_986 = {1{`RANDOM}};
  REG_986 = _RAND_986[31:0];
  _RAND_987 = {1{`RANDOM}};
  REG_987 = _RAND_987[31:0];
  _RAND_988 = {1{`RANDOM}};
  REG_988 = _RAND_988[31:0];
  _RAND_989 = {1{`RANDOM}};
  REG_989 = _RAND_989[31:0];
  _RAND_990 = {1{`RANDOM}};
  REG_990 = _RAND_990[31:0];
  _RAND_991 = {1{`RANDOM}};
  REG_991 = _RAND_991[31:0];
  _RAND_992 = {1{`RANDOM}};
  REG_992 = _RAND_992[31:0];
  _RAND_993 = {1{`RANDOM}};
  REG_993 = _RAND_993[31:0];
  _RAND_994 = {1{`RANDOM}};
  REG_994 = _RAND_994[31:0];
  _RAND_995 = {1{`RANDOM}};
  REG_995 = _RAND_995[31:0];
  _RAND_996 = {1{`RANDOM}};
  REG_996 = _RAND_996[31:0];
  _RAND_997 = {1{`RANDOM}};
  REG_997 = _RAND_997[31:0];
  _RAND_998 = {1{`RANDOM}};
  REG_998 = _RAND_998[31:0];
  _RAND_999 = {1{`RANDOM}};
  out = _RAND_999[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

